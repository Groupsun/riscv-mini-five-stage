module PC( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_addr_input, // @[:@6.4]
  input         io_pc_write, // @[:@6.4]
  output [31:0] io_pc_out // @[:@6.4]
);
  reg [31:0] PC_reg; // @[PC.scala 24:23:@8.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_14; // @[PC.scala 26:16:@10.4]
  assign _T_14 = io_pc_write ? io_addr_input : PC_reg; // @[PC.scala 26:16:@10.4]
  assign io_pc_out = PC_reg; // @[PC.scala 27:13:@12.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  PC_reg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      PC_reg <= 32'h0;
    end else begin
      if (io_pc_write) begin
        PC_reg <= io_addr_input;
      end
    end
  end
endmodule
module InstCache( // @[:@14.2]
  input         clock, // @[:@15.4]
  input  [31:0] io_addr, // @[:@17.4]
  output [31:0] io_inst // @[:@17.4]
);
  reg [7:0] cache [0:127]; // @[InstCache.scala 29:18:@19.4]
  reg [31:0] _RAND_0;
  wire [7:0] cache__T_12_data; // @[InstCache.scala 29:18:@19.4]
  wire [6:0] cache__T_12_addr; // @[InstCache.scala 29:18:@19.4]
  wire [7:0] cache__T_17_data; // @[InstCache.scala 29:18:@19.4]
  wire [6:0] cache__T_17_addr; // @[InstCache.scala 29:18:@19.4]
  wire [7:0] cache__T_22_data; // @[InstCache.scala 29:18:@19.4]
  wire [6:0] cache__T_22_addr; // @[InstCache.scala 29:18:@19.4]
  wire [7:0] cache__T_27_data; // @[InstCache.scala 29:18:@19.4]
  wire [6:0] cache__T_27_addr; // @[InstCache.scala 29:18:@19.4]
  wire [32:0] _T_14; // @[InstCache.scala 34:48:@22.4]
  wire [31:0] _T_15; // @[InstCache.scala 34:48:@23.4]
  wire [32:0] _T_19; // @[InstCache.scala 34:70:@26.4]
  wire [31:0] _T_20; // @[InstCache.scala 34:70:@27.4]
  wire [32:0] _T_24; // @[InstCache.scala 34:92:@30.4]
  wire [31:0] _T_25; // @[InstCache.scala 34:92:@31.4]
  wire [15:0] _T_28; // @[Cat.scala 30:58:@34.4]
  wire [15:0] _T_29; // @[Cat.scala 30:58:@35.4]
  assign cache__T_12_addr = io_addr[6:0];
  assign cache__T_12_data = cache[cache__T_12_addr]; // @[InstCache.scala 29:18:@19.4]
  assign cache__T_17_addr = _T_15[6:0];
  assign cache__T_17_data = cache[cache__T_17_addr]; // @[InstCache.scala 29:18:@19.4]
  assign cache__T_22_addr = _T_20[6:0];
  assign cache__T_22_data = cache[cache__T_22_addr]; // @[InstCache.scala 29:18:@19.4]
  assign cache__T_27_addr = _T_25[6:0];
  assign cache__T_27_data = cache[cache__T_27_addr]; // @[InstCache.scala 29:18:@19.4]
  assign _T_14 = io_addr + 32'h1; // @[InstCache.scala 34:48:@22.4]
  assign _T_15 = io_addr + 32'h1; // @[InstCache.scala 34:48:@23.4]
  assign _T_19 = io_addr + 32'h2; // @[InstCache.scala 34:70:@26.4]
  assign _T_20 = io_addr + 32'h2; // @[InstCache.scala 34:70:@27.4]
  assign _T_24 = io_addr + 32'h3; // @[InstCache.scala 34:92:@30.4]
  assign _T_25 = io_addr + 32'h3; // @[InstCache.scala 34:92:@31.4]
  assign _T_28 = {cache__T_22_data,cache__T_27_data}; // @[Cat.scala 30:58:@34.4]
  assign _T_29 = {cache__T_12_data,cache__T_17_data}; // @[Cat.scala 30:58:@35.4]
  assign io_inst = {_T_29,_T_28}; // @[InstCache.scala 34:11:@37.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
endmodule
module IF_ID_Register( // @[:@39.2]
  input         clock, // @[:@40.4]
  input         reset, // @[:@41.4]
  input  [31:0] io_if_pc, // @[:@42.4]
  input  [31:0] io_if_inst, // @[:@42.4]
  input         io_if_id_write, // @[:@42.4]
  input         io_if_flush, // @[:@42.4]
  input  [31:0] io_if_pc_4, // @[:@42.4]
  output [4:0]  io_id_rs1, // @[:@42.4]
  output [4:0]  io_id_rs2, // @[:@42.4]
  output [31:0] io_id_pc, // @[:@42.4]
  output [31:0] io_id_pc_4, // @[:@42.4]
  output [31:0] io_id_inst // @[:@42.4]
);
  reg [31:0] pc_reg; // @[IF_ID_Register.scala 29:26:@44.4]
  reg [31:0] _RAND_0;
  reg [31:0] inst_reg; // @[IF_ID_Register.scala 30:26:@45.4]
  reg [31:0] _RAND_1;
  reg [31:0] pc_4_reg; // @[IF_ID_Register.scala 31:26:@46.4]
  reg [31:0] _RAND_2;
  wire [31:0] _T_34; // @[IF_ID_Register.scala 34:8:@49.4]
  wire [31:0] _T_35; // @[IF_ID_Register.scala 33:16:@50.4]
  wire [31:0] _T_39; // @[IF_ID_Register.scala 37:8:@54.4]
  wire [31:0] _T_40; // @[IF_ID_Register.scala 36:18:@55.4]
  wire [31:0] _T_44; // @[IF_ID_Register.scala 40:8:@59.4]
  wire [31:0] _T_45; // @[IF_ID_Register.scala 39:18:@60.4]
  assign _T_34 = io_if_id_write ? io_if_pc : pc_reg; // @[IF_ID_Register.scala 34:8:@49.4]
  assign _T_35 = io_if_flush ? 32'h0 : _T_34; // @[IF_ID_Register.scala 33:16:@50.4]
  assign _T_39 = io_if_id_write ? io_if_inst : inst_reg; // @[IF_ID_Register.scala 37:8:@54.4]
  assign _T_40 = io_if_flush ? 32'h0 : _T_39; // @[IF_ID_Register.scala 36:18:@55.4]
  assign _T_44 = io_if_id_write ? io_if_pc_4 : pc_4_reg; // @[IF_ID_Register.scala 40:8:@59.4]
  assign _T_45 = io_if_flush ? 32'h0 : _T_44; // @[IF_ID_Register.scala 39:18:@60.4]
  assign io_id_rs1 = inst_reg[19:15]; // @[IF_ID_Register.scala 45:15:@66.4]
  assign io_id_rs2 = inst_reg[24:20]; // @[IF_ID_Register.scala 46:15:@68.4]
  assign io_id_pc = pc_reg; // @[IF_ID_Register.scala 42:15:@62.4]
  assign io_id_pc_4 = pc_4_reg; // @[IF_ID_Register.scala 43:15:@63.4]
  assign io_id_inst = inst_reg; // @[IF_ID_Register.scala 44:15:@64.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_reg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inst_reg = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  pc_4_reg = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc_reg <= 32'h0;
    end else begin
      if (io_if_flush) begin
        pc_reg <= 32'h0;
      end else begin
        if (io_if_id_write) begin
          pc_reg <= io_if_pc;
        end
      end
    end
    if (reset) begin
      inst_reg <= 32'h0;
    end else begin
      if (io_if_flush) begin
        inst_reg <= 32'h0;
      end else begin
        if (io_if_id_write) begin
          inst_reg <= io_if_inst;
        end
      end
    end
    if (reset) begin
      pc_4_reg <= 32'h0;
    end else begin
      if (io_if_flush) begin
        pc_4_reg <= 32'h0;
      end else begin
        if (io_if_id_write) begin
          pc_4_reg <= io_if_pc_4;
        end
      end
    end
  end
endmodule
module RegFile( // @[:@70.2]
  input         clock, // @[:@71.4]
  input  [4:0]  io_rs1, // @[:@73.4]
  input  [4:0]  io_rs2, // @[:@73.4]
  input  [4:0]  io_rd, // @[:@73.4]
  input  [31:0] io_wdata, // @[:@73.4]
  input         io_regwrite, // @[:@73.4]
  output [31:0] io_rs1_out, // @[:@73.4]
  output [31:0] io_rs2_out // @[:@73.4]
);
  reg [31:0] regfile [0:31]; // @[RegFile.scala 27:20:@75.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_25_data; // @[RegFile.scala 27:20:@75.4]
  wire [4:0] regfile__T_25_addr; // @[RegFile.scala 27:20:@75.4]
  wire [31:0] regfile__T_27_data; // @[RegFile.scala 27:20:@75.4]
  wire [4:0] regfile__T_27_addr; // @[RegFile.scala 27:20:@75.4]
  wire [31:0] regfile__T_34_data; // @[RegFile.scala 27:20:@75.4]
  wire [4:0] regfile__T_34_addr; // @[RegFile.scala 27:20:@75.4]
  wire [31:0] regfile__T_36_data; // @[RegFile.scala 27:20:@75.4]
  wire [4:0] regfile__T_36_addr; // @[RegFile.scala 27:20:@75.4]
  wire  regfile__T_36_mask; // @[RegFile.scala 27:20:@75.4]
  wire  regfile__T_36_en; // @[RegFile.scala 27:20:@75.4]
  wire  _T_22; // @[RegFile.scala 31:58:@77.4]
  wire  inside_forward_1; // @[RegFile.scala 31:47:@78.4]
  wire  _T_24; // @[RegFile.scala 32:58:@80.4]
  wire  inside_forward_2; // @[RegFile.scala 32:47:@81.4]
  wire  _T_31; // @[RegFile.scala 37:60:@89.4]
  wire [31:0] _T_33; // @[RegFile.scala 37:53:@90.4]
  assign regfile__T_25_addr = io_rs1;
  assign regfile__T_25_data = regfile[regfile__T_25_addr]; // @[RegFile.scala 27:20:@75.4]
  assign regfile__T_27_addr = io_rs2;
  assign regfile__T_27_data = regfile[regfile__T_27_addr]; // @[RegFile.scala 27:20:@75.4]
  assign regfile__T_34_addr = io_rd;
  assign regfile__T_34_data = regfile[regfile__T_34_addr]; // @[RegFile.scala 27:20:@75.4]
  assign regfile__T_36_data = io_regwrite ? _T_33 : regfile__T_34_data;
  assign regfile__T_36_addr = io_rd;
  assign regfile__T_36_mask = 1'h1;
  assign regfile__T_36_en = 1'h1;
  assign _T_22 = io_rs1 == io_rd; // @[RegFile.scala 31:58:@77.4]
  assign inside_forward_1 = io_regwrite & _T_22; // @[RegFile.scala 31:47:@78.4]
  assign _T_24 = io_rs2 == io_rd; // @[RegFile.scala 32:58:@80.4]
  assign inside_forward_2 = io_regwrite & _T_24; // @[RegFile.scala 32:47:@81.4]
  assign _T_31 = io_rd == 5'h0; // @[RegFile.scala 37:60:@89.4]
  assign _T_33 = _T_31 ? 32'h0 : io_wdata; // @[RegFile.scala 37:53:@90.4]
  assign io_rs1_out = inside_forward_1 ? io_wdata : regfile__T_25_data; // @[RegFile.scala 34:14:@84.4]
  assign io_rs2_out = inside_forward_2 ? io_wdata : regfile__T_27_data; // @[RegFile.scala 35:14:@87.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(regfile__T_36_en & regfile__T_36_mask) begin
      regfile[regfile__T_36_addr] <= regfile__T_36_data; // @[RegFile.scala 27:20:@75.4]
    end
  end
endmodule
module ImmGen( // @[:@96.2]
  input  [31:0] io_inst_in, // @[:@99.4]
  input  [2:0]  io_imm_sel, // @[:@99.4]
  output [31:0] io_imm // @[:@99.4]
);
  wire [11:0] _T_12; // @[ImmGen.scala 26:25:@102.4]
  wire [11:0] Iimm; // @[ImmGen.scala 26:40:@103.4]
  wire [6:0] _T_13; // @[ImmGen.scala 27:29:@104.4]
  wire [4:0] _T_14; // @[ImmGen.scala 27:49:@105.4]
  wire [11:0] _T_15; // @[Cat.scala 30:58:@106.4]
  wire [11:0] Simm; // @[ImmGen.scala 27:64:@107.4]
  wire  _T_16; // @[ImmGen.scala 28:29:@108.4]
  wire  _T_17; // @[ImmGen.scala 28:45:@109.4]
  wire [5:0] _T_18; // @[ImmGen.scala 28:60:@110.4]
  wire [3:0] _T_19; // @[ImmGen.scala 28:80:@111.4]
  wire [12:0] _T_24; // @[Cat.scala 30:58:@115.4]
  wire [12:0] SBimm; // @[ImmGen.scala 28:105:@116.4]
  wire [19:0] _T_25; // @[ImmGen.scala 29:29:@117.4]
  wire [31:0] _T_27; // @[Cat.scala 30:58:@118.4]
  wire [31:0] Uimm; // @[ImmGen.scala 29:56:@119.4]
  wire [7:0] _T_29; // @[ImmGen.scala 30:45:@121.4]
  wire  _T_30; // @[ImmGen.scala 30:65:@122.4]
  wire [9:0] _T_31; // @[ImmGen.scala 30:81:@123.4]
  wire [20:0] _T_36; // @[Cat.scala 30:58:@127.4]
  wire [20:0] UJimm; // @[ImmGen.scala 30:107:@128.4]
  wire  _T_90; // @[Mux.scala 46:19:@129.4]
  wire [20:0] _T_91; // @[Mux.scala 46:16:@130.4]
  wire  _T_92; // @[Mux.scala 46:19:@131.4]
  wire [31:0] _T_93; // @[Mux.scala 46:16:@132.4]
  wire  _T_94; // @[Mux.scala 46:19:@133.4]
  wire [31:0] _T_95; // @[Mux.scala 46:16:@134.4]
  wire  _T_96; // @[Mux.scala 46:19:@135.4]
  wire [31:0] _T_97; // @[Mux.scala 46:16:@136.4]
  wire  _T_98; // @[Mux.scala 46:19:@137.4]
  wire [31:0] _T_99; // @[Mux.scala 46:16:@138.4]
  wire  _T_100; // @[Mux.scala 46:19:@139.4]
  wire [31:0] _T_101; // @[Mux.scala 46:16:@140.4]
  assign _T_12 = io_inst_in[31:20]; // @[ImmGen.scala 26:25:@102.4]
  assign Iimm = $signed(_T_12); // @[ImmGen.scala 26:40:@103.4]
  assign _T_13 = io_inst_in[31:25]; // @[ImmGen.scala 27:29:@104.4]
  assign _T_14 = io_inst_in[11:7]; // @[ImmGen.scala 27:49:@105.4]
  assign _T_15 = {_T_13,_T_14}; // @[Cat.scala 30:58:@106.4]
  assign Simm = $signed(_T_15); // @[ImmGen.scala 27:64:@107.4]
  assign _T_16 = io_inst_in[31]; // @[ImmGen.scala 28:29:@108.4]
  assign _T_17 = io_inst_in[7]; // @[ImmGen.scala 28:45:@109.4]
  assign _T_18 = io_inst_in[30:25]; // @[ImmGen.scala 28:60:@110.4]
  assign _T_19 = io_inst_in[11:8]; // @[ImmGen.scala 28:80:@111.4]
  assign _T_24 = {_T_16,_T_17,_T_18,_T_19,1'h0}; // @[Cat.scala 30:58:@115.4]
  assign SBimm = $signed(_T_24); // @[ImmGen.scala 28:105:@116.4]
  assign _T_25 = io_inst_in[31:12]; // @[ImmGen.scala 29:29:@117.4]
  assign _T_27 = {_T_25,12'h0}; // @[Cat.scala 30:58:@118.4]
  assign Uimm = $signed(_T_27); // @[ImmGen.scala 29:56:@119.4]
  assign _T_29 = io_inst_in[19:12]; // @[ImmGen.scala 30:45:@121.4]
  assign _T_30 = io_inst_in[20]; // @[ImmGen.scala 30:65:@122.4]
  assign _T_31 = io_inst_in[30:21]; // @[ImmGen.scala 30:81:@123.4]
  assign _T_36 = {_T_16,_T_29,_T_30,_T_31,1'h0}; // @[Cat.scala 30:58:@127.4]
  assign UJimm = $signed(_T_36); // @[ImmGen.scala 30:107:@128.4]
  assign _T_90 = 3'h6 == io_imm_sel; // @[Mux.scala 46:19:@129.4]
  assign _T_91 = _T_90 ? $signed(UJimm) : $signed(21'sh0); // @[Mux.scala 46:16:@130.4]
  assign _T_92 = 3'h5 == io_imm_sel; // @[Mux.scala 46:19:@131.4]
  assign _T_93 = _T_92 ? $signed(Uimm) : $signed({{11{_T_91[20]}},_T_91}); // @[Mux.scala 46:16:@132.4]
  assign _T_94 = 3'h4 == io_imm_sel; // @[Mux.scala 46:19:@133.4]
  assign _T_95 = _T_94 ? $signed({{19{SBimm[12]}},SBimm}) : $signed(_T_93); // @[Mux.scala 46:16:@134.4]
  assign _T_96 = 3'h3 == io_imm_sel; // @[Mux.scala 46:19:@135.4]
  assign _T_97 = _T_96 ? $signed({{20{Simm[11]}},Simm}) : $signed(_T_95); // @[Mux.scala 46:16:@136.4]
  assign _T_98 = 3'h2 == io_imm_sel; // @[Mux.scala 46:19:@137.4]
  assign _T_99 = _T_98 ? $signed({{20{Iimm[11]}},Iimm}) : $signed(_T_97); // @[Mux.scala 46:16:@138.4]
  assign _T_100 = 3'h1 == io_imm_sel; // @[Mux.scala 46:19:@139.4]
  assign _T_101 = _T_100 ? $signed(32'sh0) : $signed(_T_99); // @[Mux.scala 46:16:@140.4]
  assign io_imm = $unsigned(_T_101); // @[ImmGen.scala 32:10:@142.4]
endmodule
module Control( // @[:@144.2]
  input  [31:0] io_inst, // @[:@147.4]
  output        io_Reg_Write, // @[:@147.4]
  output [2:0]  io_Imm_Sel, // @[:@147.4]
  output        io_ALU_Src, // @[:@147.4]
  output [4:0]  io_ALUOp, // @[:@147.4]
  output        io_Branch, // @[:@147.4]
  output        io_Branch_Src, // @[:@147.4]
  output        io_Mem_Read, // @[:@147.4]
  output        io_Mem_Write, // @[:@147.4]
  output [1:0]  io_Data_Size, // @[:@147.4]
  output        io_Load_Type, // @[:@147.4]
  output [2:0]  io_Mem_to_Reg, // @[:@147.4]
  output        io_Jump_Type // @[:@147.4]
);
  wire [31:0] _T_33; // @[Lookup.scala 9:38:@149.4]
  wire  _T_34; // @[Lookup.scala 9:38:@150.4]
  wire  _T_38; // @[Lookup.scala 9:38:@152.4]
  wire  _T_42; // @[Lookup.scala 9:38:@154.4]
  wire  _T_46; // @[Lookup.scala 9:38:@156.4]
  wire  _T_50; // @[Lookup.scala 9:38:@158.4]
  wire [31:0] _T_53; // @[Lookup.scala 9:38:@159.4]
  wire  _T_54; // @[Lookup.scala 9:38:@160.4]
  wire  _T_58; // @[Lookup.scala 9:38:@162.4]
  wire  _T_62; // @[Lookup.scala 9:38:@164.4]
  wire  _T_66; // @[Lookup.scala 9:38:@166.4]
  wire  _T_70; // @[Lookup.scala 9:38:@168.4]
  wire  _T_74; // @[Lookup.scala 9:38:@170.4]
  wire  _T_78; // @[Lookup.scala 9:38:@172.4]
  wire  _T_82; // @[Lookup.scala 9:38:@174.4]
  wire  _T_86; // @[Lookup.scala 9:38:@176.4]
  wire  _T_90; // @[Lookup.scala 9:38:@178.4]
  wire  _T_94; // @[Lookup.scala 9:38:@180.4]
  wire  _T_98; // @[Lookup.scala 9:38:@182.4]
  wire  _T_102; // @[Lookup.scala 9:38:@184.4]
  wire  _T_106; // @[Lookup.scala 9:38:@186.4]
  wire  _T_110; // @[Lookup.scala 9:38:@188.4]
  wire  _T_114; // @[Lookup.scala 9:38:@190.4]
  wire  _T_118; // @[Lookup.scala 9:38:@192.4]
  wire  _T_122; // @[Lookup.scala 9:38:@194.4]
  wire  _T_126; // @[Lookup.scala 9:38:@196.4]
  wire  _T_130; // @[Lookup.scala 9:38:@198.4]
  wire  _T_134; // @[Lookup.scala 9:38:@200.4]
  wire  _T_138; // @[Lookup.scala 9:38:@202.4]
  wire  _T_142; // @[Lookup.scala 9:38:@204.4]
  wire  _T_146; // @[Lookup.scala 9:38:@206.4]
  wire  _T_150; // @[Lookup.scala 9:38:@208.4]
  wire  _T_154; // @[Lookup.scala 9:38:@210.4]
  wire  _T_158; // @[Lookup.scala 9:38:@212.4]
  wire  _T_162; // @[Lookup.scala 9:38:@214.4]
  wire [31:0] _T_165; // @[Lookup.scala 9:38:@215.4]
  wire  _T_166; // @[Lookup.scala 9:38:@216.4]
  wire  _T_170; // @[Lookup.scala 9:38:@218.4]
  wire  _T_174; // @[Lookup.scala 9:38:@220.4]
  wire  _T_178; // @[Lookup.scala 9:38:@222.4]
  wire  _T_185; // @[Lookup.scala 11:37:@227.4]
  wire  _T_186; // @[Lookup.scala 11:37:@228.4]
  wire  _T_187; // @[Lookup.scala 11:37:@229.4]
  wire  _T_188; // @[Lookup.scala 11:37:@230.4]
  wire  _T_189; // @[Lookup.scala 11:37:@231.4]
  wire  _T_190; // @[Lookup.scala 11:37:@232.4]
  wire  _T_191; // @[Lookup.scala 11:37:@233.4]
  wire  _T_192; // @[Lookup.scala 11:37:@234.4]
  wire  _T_193; // @[Lookup.scala 11:37:@235.4]
  wire  _T_194; // @[Lookup.scala 11:37:@236.4]
  wire  _T_195; // @[Lookup.scala 11:37:@237.4]
  wire  _T_196; // @[Lookup.scala 11:37:@238.4]
  wire  _T_197; // @[Lookup.scala 11:37:@239.4]
  wire  _T_198; // @[Lookup.scala 11:37:@240.4]
  wire  _T_199; // @[Lookup.scala 11:37:@241.4]
  wire  _T_200; // @[Lookup.scala 11:37:@242.4]
  wire  _T_201; // @[Lookup.scala 11:37:@243.4]
  wire  _T_202; // @[Lookup.scala 11:37:@244.4]
  wire  _T_203; // @[Lookup.scala 11:37:@245.4]
  wire  _T_204; // @[Lookup.scala 11:37:@246.4]
  wire  _T_205; // @[Lookup.scala 11:37:@247.4]
  wire  _T_206; // @[Lookup.scala 11:37:@248.4]
  wire  _T_207; // @[Lookup.scala 11:37:@249.4]
  wire  _T_208; // @[Lookup.scala 11:37:@250.4]
  wire  _T_209; // @[Lookup.scala 11:37:@251.4]
  wire  _T_210; // @[Lookup.scala 11:37:@252.4]
  wire  _T_211; // @[Lookup.scala 11:37:@253.4]
  wire  _T_212; // @[Lookup.scala 11:37:@254.4]
  wire  _T_213; // @[Lookup.scala 11:37:@255.4]
  wire  _T_214; // @[Lookup.scala 11:37:@256.4]
  wire  _T_215; // @[Lookup.scala 11:37:@257.4]
  wire  _T_216; // @[Lookup.scala 11:37:@258.4]
  wire  _T_217; // @[Lookup.scala 11:37:@259.4]
  wire  _T_218; // @[Lookup.scala 11:37:@260.4]
  wire  _T_219; // @[Lookup.scala 11:37:@261.4]
  wire [2:0] _T_221; // @[Lookup.scala 11:37:@264.4]
  wire [2:0] _T_222; // @[Lookup.scala 11:37:@265.4]
  wire [2:0] _T_223; // @[Lookup.scala 11:37:@266.4]
  wire [2:0] _T_224; // @[Lookup.scala 11:37:@267.4]
  wire [2:0] _T_225; // @[Lookup.scala 11:37:@268.4]
  wire [2:0] _T_226; // @[Lookup.scala 11:37:@269.4]
  wire [2:0] _T_227; // @[Lookup.scala 11:37:@270.4]
  wire [2:0] _T_228; // @[Lookup.scala 11:37:@271.4]
  wire [2:0] _T_229; // @[Lookup.scala 11:37:@272.4]
  wire [2:0] _T_230; // @[Lookup.scala 11:37:@273.4]
  wire [2:0] _T_231; // @[Lookup.scala 11:37:@274.4]
  wire [2:0] _T_232; // @[Lookup.scala 11:37:@275.4]
  wire [2:0] _T_233; // @[Lookup.scala 11:37:@276.4]
  wire [2:0] _T_234; // @[Lookup.scala 11:37:@277.4]
  wire [2:0] _T_235; // @[Lookup.scala 11:37:@278.4]
  wire [2:0] _T_236; // @[Lookup.scala 11:37:@279.4]
  wire [2:0] _T_237; // @[Lookup.scala 11:37:@280.4]
  wire [2:0] _T_238; // @[Lookup.scala 11:37:@281.4]
  wire [2:0] _T_239; // @[Lookup.scala 11:37:@282.4]
  wire [2:0] _T_240; // @[Lookup.scala 11:37:@283.4]
  wire [2:0] _T_241; // @[Lookup.scala 11:37:@284.4]
  wire [2:0] _T_242; // @[Lookup.scala 11:37:@285.4]
  wire [2:0] _T_243; // @[Lookup.scala 11:37:@286.4]
  wire [2:0] _T_244; // @[Lookup.scala 11:37:@287.4]
  wire [2:0] _T_245; // @[Lookup.scala 11:37:@288.4]
  wire [2:0] _T_246; // @[Lookup.scala 11:37:@289.4]
  wire [2:0] _T_247; // @[Lookup.scala 11:37:@290.4]
  wire [2:0] _T_248; // @[Lookup.scala 11:37:@291.4]
  wire [2:0] _T_249; // @[Lookup.scala 11:37:@292.4]
  wire [2:0] _T_250; // @[Lookup.scala 11:37:@293.4]
  wire [2:0] _T_251; // @[Lookup.scala 11:37:@294.4]
  wire [2:0] _T_252; // @[Lookup.scala 11:37:@295.4]
  wire [2:0] _T_253; // @[Lookup.scala 11:37:@296.4]
  wire [2:0] _T_254; // @[Lookup.scala 11:37:@297.4]
  wire [2:0] _T_255; // @[Lookup.scala 11:37:@298.4]
  wire [2:0] _T_256; // @[Lookup.scala 11:37:@299.4]
  wire  _T_269; // @[Lookup.scala 11:37:@313.4]
  wire  _T_270; // @[Lookup.scala 11:37:@314.4]
  wire  _T_271; // @[Lookup.scala 11:37:@315.4]
  wire  _T_272; // @[Lookup.scala 11:37:@316.4]
  wire  _T_273; // @[Lookup.scala 11:37:@317.4]
  wire  _T_274; // @[Lookup.scala 11:37:@318.4]
  wire  _T_275; // @[Lookup.scala 11:37:@319.4]
  wire  _T_276; // @[Lookup.scala 11:37:@320.4]
  wire  _T_277; // @[Lookup.scala 11:37:@321.4]
  wire  _T_278; // @[Lookup.scala 11:37:@322.4]
  wire  _T_279; // @[Lookup.scala 11:37:@323.4]
  wire  _T_280; // @[Lookup.scala 11:37:@324.4]
  wire  _T_281; // @[Lookup.scala 11:37:@325.4]
  wire  _T_282; // @[Lookup.scala 11:37:@326.4]
  wire  _T_283; // @[Lookup.scala 11:37:@327.4]
  wire  _T_284; // @[Lookup.scala 11:37:@328.4]
  wire  _T_285; // @[Lookup.scala 11:37:@329.4]
  wire  _T_286; // @[Lookup.scala 11:37:@330.4]
  wire  _T_287; // @[Lookup.scala 11:37:@331.4]
  wire  _T_288; // @[Lookup.scala 11:37:@332.4]
  wire  _T_289; // @[Lookup.scala 11:37:@333.4]
  wire  _T_290; // @[Lookup.scala 11:37:@334.4]
  wire  _T_291; // @[Lookup.scala 11:37:@335.4]
  wire  _T_292; // @[Lookup.scala 11:37:@336.4]
  wire  _T_293; // @[Lookup.scala 11:37:@337.4]
  wire [4:0] _T_295; // @[Lookup.scala 11:37:@340.4]
  wire [4:0] _T_296; // @[Lookup.scala 11:37:@341.4]
  wire [4:0] _T_297; // @[Lookup.scala 11:37:@342.4]
  wire [4:0] _T_298; // @[Lookup.scala 11:37:@343.4]
  wire [4:0] _T_299; // @[Lookup.scala 11:37:@344.4]
  wire [4:0] _T_300; // @[Lookup.scala 11:37:@345.4]
  wire [4:0] _T_301; // @[Lookup.scala 11:37:@346.4]
  wire [4:0] _T_302; // @[Lookup.scala 11:37:@347.4]
  wire [4:0] _T_303; // @[Lookup.scala 11:37:@348.4]
  wire [4:0] _T_304; // @[Lookup.scala 11:37:@349.4]
  wire [4:0] _T_305; // @[Lookup.scala 11:37:@350.4]
  wire [4:0] _T_306; // @[Lookup.scala 11:37:@351.4]
  wire [4:0] _T_307; // @[Lookup.scala 11:37:@352.4]
  wire [4:0] _T_308; // @[Lookup.scala 11:37:@353.4]
  wire [4:0] _T_309; // @[Lookup.scala 11:37:@354.4]
  wire [4:0] _T_310; // @[Lookup.scala 11:37:@355.4]
  wire [4:0] _T_311; // @[Lookup.scala 11:37:@356.4]
  wire [4:0] _T_312; // @[Lookup.scala 11:37:@357.4]
  wire [4:0] _T_313; // @[Lookup.scala 11:37:@358.4]
  wire [4:0] _T_314; // @[Lookup.scala 11:37:@359.4]
  wire [4:0] _T_315; // @[Lookup.scala 11:37:@360.4]
  wire [4:0] _T_316; // @[Lookup.scala 11:37:@361.4]
  wire [4:0] _T_317; // @[Lookup.scala 11:37:@362.4]
  wire [4:0] _T_318; // @[Lookup.scala 11:37:@363.4]
  wire [4:0] _T_319; // @[Lookup.scala 11:37:@364.4]
  wire [4:0] _T_320; // @[Lookup.scala 11:37:@365.4]
  wire [4:0] _T_321; // @[Lookup.scala 11:37:@366.4]
  wire [4:0] _T_322; // @[Lookup.scala 11:37:@367.4]
  wire [4:0] _T_323; // @[Lookup.scala 11:37:@368.4]
  wire [4:0] _T_324; // @[Lookup.scala 11:37:@369.4]
  wire [4:0] _T_325; // @[Lookup.scala 11:37:@370.4]
  wire [4:0] _T_326; // @[Lookup.scala 11:37:@371.4]
  wire [4:0] _T_327; // @[Lookup.scala 11:37:@372.4]
  wire [4:0] _T_328; // @[Lookup.scala 11:37:@373.4]
  wire [4:0] _T_329; // @[Lookup.scala 11:37:@374.4]
  wire [4:0] _T_330; // @[Lookup.scala 11:37:@375.4]
  wire  _T_335; // @[Lookup.scala 11:37:@381.4]
  wire  _T_336; // @[Lookup.scala 11:37:@382.4]
  wire  _T_337; // @[Lookup.scala 11:37:@383.4]
  wire  _T_338; // @[Lookup.scala 11:37:@384.4]
  wire  _T_339; // @[Lookup.scala 11:37:@385.4]
  wire  _T_340; // @[Lookup.scala 11:37:@386.4]
  wire  _T_341; // @[Lookup.scala 11:37:@387.4]
  wire  _T_342; // @[Lookup.scala 11:37:@388.4]
  wire  _T_343; // @[Lookup.scala 11:37:@389.4]
  wire  _T_344; // @[Lookup.scala 11:37:@390.4]
  wire  _T_345; // @[Lookup.scala 11:37:@391.4]
  wire  _T_346; // @[Lookup.scala 11:37:@392.4]
  wire  _T_347; // @[Lookup.scala 11:37:@393.4]
  wire  _T_348; // @[Lookup.scala 11:37:@394.4]
  wire  _T_349; // @[Lookup.scala 11:37:@395.4]
  wire  _T_350; // @[Lookup.scala 11:37:@396.4]
  wire  _T_351; // @[Lookup.scala 11:37:@397.4]
  wire  _T_352; // @[Lookup.scala 11:37:@398.4]
  wire  _T_353; // @[Lookup.scala 11:37:@399.4]
  wire  _T_354; // @[Lookup.scala 11:37:@400.4]
  wire  _T_355; // @[Lookup.scala 11:37:@401.4]
  wire  _T_356; // @[Lookup.scala 11:37:@402.4]
  wire  _T_357; // @[Lookup.scala 11:37:@403.4]
  wire  _T_358; // @[Lookup.scala 11:37:@404.4]
  wire  _T_359; // @[Lookup.scala 11:37:@405.4]
  wire  _T_360; // @[Lookup.scala 11:37:@406.4]
  wire  _T_361; // @[Lookup.scala 11:37:@407.4]
  wire  _T_362; // @[Lookup.scala 11:37:@408.4]
  wire  _T_363; // @[Lookup.scala 11:37:@409.4]
  wire  _T_364; // @[Lookup.scala 11:37:@410.4]
  wire  _T_365; // @[Lookup.scala 11:37:@411.4]
  wire  _T_366; // @[Lookup.scala 11:37:@412.4]
  wire  _T_367; // @[Lookup.scala 11:37:@413.4]
  wire  _T_372; // @[Lookup.scala 11:37:@419.4]
  wire  _T_373; // @[Lookup.scala 11:37:@420.4]
  wire  _T_374; // @[Lookup.scala 11:37:@421.4]
  wire  _T_375; // @[Lookup.scala 11:37:@422.4]
  wire  _T_376; // @[Lookup.scala 11:37:@423.4]
  wire  _T_377; // @[Lookup.scala 11:37:@424.4]
  wire  _T_378; // @[Lookup.scala 11:37:@425.4]
  wire  _T_379; // @[Lookup.scala 11:37:@426.4]
  wire  _T_380; // @[Lookup.scala 11:37:@427.4]
  wire  _T_381; // @[Lookup.scala 11:37:@428.4]
  wire  _T_382; // @[Lookup.scala 11:37:@429.4]
  wire  _T_383; // @[Lookup.scala 11:37:@430.4]
  wire  _T_384; // @[Lookup.scala 11:37:@431.4]
  wire  _T_385; // @[Lookup.scala 11:37:@432.4]
  wire  _T_386; // @[Lookup.scala 11:37:@433.4]
  wire  _T_387; // @[Lookup.scala 11:37:@434.4]
  wire  _T_388; // @[Lookup.scala 11:37:@435.4]
  wire  _T_389; // @[Lookup.scala 11:37:@436.4]
  wire  _T_390; // @[Lookup.scala 11:37:@437.4]
  wire  _T_391; // @[Lookup.scala 11:37:@438.4]
  wire  _T_392; // @[Lookup.scala 11:37:@439.4]
  wire  _T_393; // @[Lookup.scala 11:37:@440.4]
  wire  _T_394; // @[Lookup.scala 11:37:@441.4]
  wire  _T_395; // @[Lookup.scala 11:37:@442.4]
  wire  _T_396; // @[Lookup.scala 11:37:@443.4]
  wire  _T_397; // @[Lookup.scala 11:37:@444.4]
  wire  _T_398; // @[Lookup.scala 11:37:@445.4]
  wire  _T_399; // @[Lookup.scala 11:37:@446.4]
  wire  _T_400; // @[Lookup.scala 11:37:@447.4]
  wire  _T_401; // @[Lookup.scala 11:37:@448.4]
  wire  _T_402; // @[Lookup.scala 11:37:@449.4]
  wire  _T_403; // @[Lookup.scala 11:37:@450.4]
  wire  _T_404; // @[Lookup.scala 11:37:@451.4]
  wire  _T_420; // @[Lookup.scala 11:37:@468.4]
  wire  _T_421; // @[Lookup.scala 11:37:@469.4]
  wire  _T_422; // @[Lookup.scala 11:37:@470.4]
  wire  _T_423; // @[Lookup.scala 11:37:@471.4]
  wire  _T_424; // @[Lookup.scala 11:37:@472.4]
  wire  _T_425; // @[Lookup.scala 11:37:@473.4]
  wire  _T_426; // @[Lookup.scala 11:37:@474.4]
  wire  _T_427; // @[Lookup.scala 11:37:@475.4]
  wire  _T_428; // @[Lookup.scala 11:37:@476.4]
  wire  _T_429; // @[Lookup.scala 11:37:@477.4]
  wire  _T_430; // @[Lookup.scala 11:37:@478.4]
  wire  _T_431; // @[Lookup.scala 11:37:@479.4]
  wire  _T_432; // @[Lookup.scala 11:37:@480.4]
  wire  _T_433; // @[Lookup.scala 11:37:@481.4]
  wire  _T_434; // @[Lookup.scala 11:37:@482.4]
  wire  _T_435; // @[Lookup.scala 11:37:@483.4]
  wire  _T_436; // @[Lookup.scala 11:37:@484.4]
  wire  _T_437; // @[Lookup.scala 11:37:@485.4]
  wire  _T_438; // @[Lookup.scala 11:37:@486.4]
  wire  _T_439; // @[Lookup.scala 11:37:@487.4]
  wire  _T_440; // @[Lookup.scala 11:37:@488.4]
  wire  _T_441; // @[Lookup.scala 11:37:@489.4]
  wire  _T_456; // @[Lookup.scala 11:37:@505.4]
  wire  _T_457; // @[Lookup.scala 11:37:@506.4]
  wire  _T_458; // @[Lookup.scala 11:37:@507.4]
  wire  _T_459; // @[Lookup.scala 11:37:@508.4]
  wire  _T_460; // @[Lookup.scala 11:37:@509.4]
  wire  _T_461; // @[Lookup.scala 11:37:@510.4]
  wire  _T_462; // @[Lookup.scala 11:37:@511.4]
  wire  _T_463; // @[Lookup.scala 11:37:@512.4]
  wire  _T_464; // @[Lookup.scala 11:37:@513.4]
  wire  _T_465; // @[Lookup.scala 11:37:@514.4]
  wire  _T_466; // @[Lookup.scala 11:37:@515.4]
  wire  _T_467; // @[Lookup.scala 11:37:@516.4]
  wire  _T_468; // @[Lookup.scala 11:37:@517.4]
  wire  _T_469; // @[Lookup.scala 11:37:@518.4]
  wire  _T_470; // @[Lookup.scala 11:37:@519.4]
  wire  _T_471; // @[Lookup.scala 11:37:@520.4]
  wire  _T_472; // @[Lookup.scala 11:37:@521.4]
  wire  _T_473; // @[Lookup.scala 11:37:@522.4]
  wire  _T_474; // @[Lookup.scala 11:37:@523.4]
  wire  _T_475; // @[Lookup.scala 11:37:@524.4]
  wire  _T_476; // @[Lookup.scala 11:37:@525.4]
  wire  _T_477; // @[Lookup.scala 11:37:@526.4]
  wire  _T_478; // @[Lookup.scala 11:37:@527.4]
  wire [1:0] _T_490; // @[Lookup.scala 11:37:@540.4]
  wire [1:0] _T_491; // @[Lookup.scala 11:37:@541.4]
  wire [1:0] _T_492; // @[Lookup.scala 11:37:@542.4]
  wire [1:0] _T_493; // @[Lookup.scala 11:37:@543.4]
  wire [1:0] _T_494; // @[Lookup.scala 11:37:@544.4]
  wire [1:0] _T_495; // @[Lookup.scala 11:37:@545.4]
  wire [1:0] _T_496; // @[Lookup.scala 11:37:@546.4]
  wire [1:0] _T_497; // @[Lookup.scala 11:37:@547.4]
  wire [1:0] _T_498; // @[Lookup.scala 11:37:@548.4]
  wire [1:0] _T_499; // @[Lookup.scala 11:37:@549.4]
  wire [1:0] _T_500; // @[Lookup.scala 11:37:@550.4]
  wire [1:0] _T_501; // @[Lookup.scala 11:37:@551.4]
  wire [1:0] _T_502; // @[Lookup.scala 11:37:@552.4]
  wire [1:0] _T_503; // @[Lookup.scala 11:37:@553.4]
  wire [1:0] _T_504; // @[Lookup.scala 11:37:@554.4]
  wire [1:0] _T_505; // @[Lookup.scala 11:37:@555.4]
  wire [1:0] _T_506; // @[Lookup.scala 11:37:@556.4]
  wire [1:0] _T_507; // @[Lookup.scala 11:37:@557.4]
  wire [1:0] _T_508; // @[Lookup.scala 11:37:@558.4]
  wire [1:0] _T_509; // @[Lookup.scala 11:37:@559.4]
  wire [1:0] _T_510; // @[Lookup.scala 11:37:@560.4]
  wire [1:0] _T_511; // @[Lookup.scala 11:37:@561.4]
  wire [1:0] _T_512; // @[Lookup.scala 11:37:@562.4]
  wire [1:0] _T_513; // @[Lookup.scala 11:37:@563.4]
  wire [1:0] _T_514; // @[Lookup.scala 11:37:@564.4]
  wire [1:0] _T_515; // @[Lookup.scala 11:37:@565.4]
  wire  _T_532; // @[Lookup.scala 11:37:@583.4]
  wire  _T_533; // @[Lookup.scala 11:37:@584.4]
  wire  _T_534; // @[Lookup.scala 11:37:@585.4]
  wire  _T_535; // @[Lookup.scala 11:37:@586.4]
  wire  _T_536; // @[Lookup.scala 11:37:@587.4]
  wire  _T_537; // @[Lookup.scala 11:37:@588.4]
  wire  _T_538; // @[Lookup.scala 11:37:@589.4]
  wire  _T_539; // @[Lookup.scala 11:37:@590.4]
  wire  _T_540; // @[Lookup.scala 11:37:@591.4]
  wire  _T_541; // @[Lookup.scala 11:37:@592.4]
  wire  _T_542; // @[Lookup.scala 11:37:@593.4]
  wire  _T_543; // @[Lookup.scala 11:37:@594.4]
  wire  _T_544; // @[Lookup.scala 11:37:@595.4]
  wire  _T_545; // @[Lookup.scala 11:37:@596.4]
  wire  _T_546; // @[Lookup.scala 11:37:@597.4]
  wire  _T_547; // @[Lookup.scala 11:37:@598.4]
  wire  _T_548; // @[Lookup.scala 11:37:@599.4]
  wire  _T_549; // @[Lookup.scala 11:37:@600.4]
  wire  _T_550; // @[Lookup.scala 11:37:@601.4]
  wire  _T_551; // @[Lookup.scala 11:37:@602.4]
  wire  _T_552; // @[Lookup.scala 11:37:@603.4]
  wire [2:0] _T_554; // @[Lookup.scala 11:37:@606.4]
  wire [2:0] _T_555; // @[Lookup.scala 11:37:@607.4]
  wire [2:0] _T_556; // @[Lookup.scala 11:37:@608.4]
  wire [2:0] _T_557; // @[Lookup.scala 11:37:@609.4]
  wire [2:0] _T_558; // @[Lookup.scala 11:37:@610.4]
  wire [2:0] _T_559; // @[Lookup.scala 11:37:@611.4]
  wire [2:0] _T_560; // @[Lookup.scala 11:37:@612.4]
  wire [2:0] _T_561; // @[Lookup.scala 11:37:@613.4]
  wire [2:0] _T_562; // @[Lookup.scala 11:37:@614.4]
  wire [2:0] _T_563; // @[Lookup.scala 11:37:@615.4]
  wire [2:0] _T_564; // @[Lookup.scala 11:37:@616.4]
  wire [2:0] _T_565; // @[Lookup.scala 11:37:@617.4]
  wire [2:0] _T_566; // @[Lookup.scala 11:37:@618.4]
  wire [2:0] _T_567; // @[Lookup.scala 11:37:@619.4]
  wire [2:0] _T_568; // @[Lookup.scala 11:37:@620.4]
  wire [2:0] _T_569; // @[Lookup.scala 11:37:@621.4]
  wire [2:0] _T_570; // @[Lookup.scala 11:37:@622.4]
  wire [2:0] _T_571; // @[Lookup.scala 11:37:@623.4]
  wire [2:0] _T_572; // @[Lookup.scala 11:37:@624.4]
  wire [2:0] _T_573; // @[Lookup.scala 11:37:@625.4]
  wire [2:0] _T_574; // @[Lookup.scala 11:37:@626.4]
  wire [2:0] _T_575; // @[Lookup.scala 11:37:@627.4]
  wire [2:0] _T_576; // @[Lookup.scala 11:37:@628.4]
  wire [2:0] _T_577; // @[Lookup.scala 11:37:@629.4]
  wire [2:0] _T_578; // @[Lookup.scala 11:37:@630.4]
  wire [2:0] _T_579; // @[Lookup.scala 11:37:@631.4]
  wire [2:0] _T_580; // @[Lookup.scala 11:37:@632.4]
  wire [2:0] _T_581; // @[Lookup.scala 11:37:@633.4]
  wire [2:0] _T_582; // @[Lookup.scala 11:37:@634.4]
  wire [2:0] _T_583; // @[Lookup.scala 11:37:@635.4]
  wire [2:0] _T_584; // @[Lookup.scala 11:37:@636.4]
  wire [2:0] _T_585; // @[Lookup.scala 11:37:@637.4]
  wire [2:0] _T_586; // @[Lookup.scala 11:37:@638.4]
  wire [2:0] _T_587; // @[Lookup.scala 11:37:@639.4]
  wire [2:0] _T_588; // @[Lookup.scala 11:37:@640.4]
  wire [2:0] _T_589; // @[Lookup.scala 11:37:@641.4]
  wire  _T_595; // @[Lookup.scala 11:37:@648.4]
  wire  _T_596; // @[Lookup.scala 11:37:@649.4]
  wire  _T_597; // @[Lookup.scala 11:37:@650.4]
  wire  _T_598; // @[Lookup.scala 11:37:@651.4]
  wire  _T_599; // @[Lookup.scala 11:37:@652.4]
  wire  _T_600; // @[Lookup.scala 11:37:@653.4]
  wire  _T_601; // @[Lookup.scala 11:37:@654.4]
  wire  _T_602; // @[Lookup.scala 11:37:@655.4]
  wire  _T_603; // @[Lookup.scala 11:37:@656.4]
  wire  _T_604; // @[Lookup.scala 11:37:@657.4]
  wire  _T_605; // @[Lookup.scala 11:37:@658.4]
  wire  _T_606; // @[Lookup.scala 11:37:@659.4]
  wire  _T_607; // @[Lookup.scala 11:37:@660.4]
  wire  _T_608; // @[Lookup.scala 11:37:@661.4]
  wire  _T_609; // @[Lookup.scala 11:37:@662.4]
  wire  _T_610; // @[Lookup.scala 11:37:@663.4]
  wire  _T_611; // @[Lookup.scala 11:37:@664.4]
  wire  _T_612; // @[Lookup.scala 11:37:@665.4]
  wire  _T_613; // @[Lookup.scala 11:37:@666.4]
  wire  _T_614; // @[Lookup.scala 11:37:@667.4]
  wire  _T_615; // @[Lookup.scala 11:37:@668.4]
  wire  _T_616; // @[Lookup.scala 11:37:@669.4]
  wire  _T_617; // @[Lookup.scala 11:37:@670.4]
  wire  _T_618; // @[Lookup.scala 11:37:@671.4]
  wire  _T_619; // @[Lookup.scala 11:37:@672.4]
  wire  _T_620; // @[Lookup.scala 11:37:@673.4]
  wire  _T_621; // @[Lookup.scala 11:37:@674.4]
  wire  _T_622; // @[Lookup.scala 11:37:@675.4]
  wire  _T_623; // @[Lookup.scala 11:37:@676.4]
  wire  _T_624; // @[Lookup.scala 11:37:@677.4]
  wire  _T_625; // @[Lookup.scala 11:37:@678.4]
  wire  _T_626; // @[Lookup.scala 11:37:@679.4]
  assign _T_33 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@149.4]
  assign _T_34 = 32'h33 == _T_33; // @[Lookup.scala 9:38:@150.4]
  assign _T_38 = 32'h40000033 == _T_33; // @[Lookup.scala 9:38:@152.4]
  assign _T_42 = 32'h7033 == _T_33; // @[Lookup.scala 9:38:@154.4]
  assign _T_46 = 32'h6033 == _T_33; // @[Lookup.scala 9:38:@156.4]
  assign _T_50 = 32'h4033 == _T_33; // @[Lookup.scala 9:38:@158.4]
  assign _T_53 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@159.4]
  assign _T_54 = 32'h13 == _T_53; // @[Lookup.scala 9:38:@160.4]
  assign _T_58 = 32'h7013 == _T_53; // @[Lookup.scala 9:38:@162.4]
  assign _T_62 = 32'h6013 == _T_53; // @[Lookup.scala 9:38:@164.4]
  assign _T_66 = 32'h4013 == _T_53; // @[Lookup.scala 9:38:@166.4]
  assign _T_70 = 32'h1033 == _T_33; // @[Lookup.scala 9:38:@168.4]
  assign _T_74 = 32'h5033 == _T_33; // @[Lookup.scala 9:38:@170.4]
  assign _T_78 = 32'h40005033 == _T_33; // @[Lookup.scala 9:38:@172.4]
  assign _T_82 = 32'h1013 == _T_33; // @[Lookup.scala 9:38:@174.4]
  assign _T_86 = 32'h5013 == _T_33; // @[Lookup.scala 9:38:@176.4]
  assign _T_90 = 32'h40005013 == _T_33; // @[Lookup.scala 9:38:@178.4]
  assign _T_94 = 32'h2033 == _T_33; // @[Lookup.scala 9:38:@180.4]
  assign _T_98 = 32'h3033 == _T_33; // @[Lookup.scala 9:38:@182.4]
  assign _T_102 = 32'h2013 == _T_53; // @[Lookup.scala 9:38:@184.4]
  assign _T_106 = 32'h3013 == _T_53; // @[Lookup.scala 9:38:@186.4]
  assign _T_110 = 32'h2003 == _T_53; // @[Lookup.scala 9:38:@188.4]
  assign _T_114 = 32'h1003 == _T_53; // @[Lookup.scala 9:38:@190.4]
  assign _T_118 = 32'h3 == _T_53; // @[Lookup.scala 9:38:@192.4]
  assign _T_122 = 32'h5003 == _T_53; // @[Lookup.scala 9:38:@194.4]
  assign _T_126 = 32'h4003 == _T_53; // @[Lookup.scala 9:38:@196.4]
  assign _T_130 = 32'h2023 == _T_53; // @[Lookup.scala 9:38:@198.4]
  assign _T_134 = 32'h1023 == _T_53; // @[Lookup.scala 9:38:@200.4]
  assign _T_138 = 32'h23 == _T_53; // @[Lookup.scala 9:38:@202.4]
  assign _T_142 = 32'h63 == _T_53; // @[Lookup.scala 9:38:@204.4]
  assign _T_146 = 32'h1063 == _T_53; // @[Lookup.scala 9:38:@206.4]
  assign _T_150 = 32'h4063 == _T_53; // @[Lookup.scala 9:38:@208.4]
  assign _T_154 = 32'h5063 == _T_53; // @[Lookup.scala 9:38:@210.4]
  assign _T_158 = 32'h6063 == _T_53; // @[Lookup.scala 9:38:@212.4]
  assign _T_162 = 32'h7063 == _T_53; // @[Lookup.scala 9:38:@214.4]
  assign _T_165 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@215.4]
  assign _T_166 = 32'h6f == _T_165; // @[Lookup.scala 9:38:@216.4]
  assign _T_170 = 32'h67 == _T_53; // @[Lookup.scala 9:38:@218.4]
  assign _T_174 = 32'h37 == _T_165; // @[Lookup.scala 9:38:@220.4]
  assign _T_178 = 32'h17 == _T_165; // @[Lookup.scala 9:38:@222.4]
  assign _T_185 = _T_174 ? 1'h1 : _T_178; // @[Lookup.scala 11:37:@227.4]
  assign _T_186 = _T_170 ? 1'h1 : _T_185; // @[Lookup.scala 11:37:@228.4]
  assign _T_187 = _T_166 ? 1'h1 : _T_186; // @[Lookup.scala 11:37:@229.4]
  assign _T_188 = _T_162 ? 1'h0 : _T_187; // @[Lookup.scala 11:37:@230.4]
  assign _T_189 = _T_158 ? 1'h0 : _T_188; // @[Lookup.scala 11:37:@231.4]
  assign _T_190 = _T_154 ? 1'h0 : _T_189; // @[Lookup.scala 11:37:@232.4]
  assign _T_191 = _T_150 ? 1'h0 : _T_190; // @[Lookup.scala 11:37:@233.4]
  assign _T_192 = _T_146 ? 1'h0 : _T_191; // @[Lookup.scala 11:37:@234.4]
  assign _T_193 = _T_142 ? 1'h0 : _T_192; // @[Lookup.scala 11:37:@235.4]
  assign _T_194 = _T_138 ? 1'h0 : _T_193; // @[Lookup.scala 11:37:@236.4]
  assign _T_195 = _T_134 ? 1'h0 : _T_194; // @[Lookup.scala 11:37:@237.4]
  assign _T_196 = _T_130 ? 1'h0 : _T_195; // @[Lookup.scala 11:37:@238.4]
  assign _T_197 = _T_126 ? 1'h1 : _T_196; // @[Lookup.scala 11:37:@239.4]
  assign _T_198 = _T_122 ? 1'h1 : _T_197; // @[Lookup.scala 11:37:@240.4]
  assign _T_199 = _T_118 ? 1'h1 : _T_198; // @[Lookup.scala 11:37:@241.4]
  assign _T_200 = _T_114 ? 1'h1 : _T_199; // @[Lookup.scala 11:37:@242.4]
  assign _T_201 = _T_110 ? 1'h1 : _T_200; // @[Lookup.scala 11:37:@243.4]
  assign _T_202 = _T_106 ? 1'h1 : _T_201; // @[Lookup.scala 11:37:@244.4]
  assign _T_203 = _T_102 ? 1'h1 : _T_202; // @[Lookup.scala 11:37:@245.4]
  assign _T_204 = _T_98 ? 1'h1 : _T_203; // @[Lookup.scala 11:37:@246.4]
  assign _T_205 = _T_94 ? 1'h1 : _T_204; // @[Lookup.scala 11:37:@247.4]
  assign _T_206 = _T_90 ? 1'h1 : _T_205; // @[Lookup.scala 11:37:@248.4]
  assign _T_207 = _T_86 ? 1'h1 : _T_206; // @[Lookup.scala 11:37:@249.4]
  assign _T_208 = _T_82 ? 1'h1 : _T_207; // @[Lookup.scala 11:37:@250.4]
  assign _T_209 = _T_78 ? 1'h1 : _T_208; // @[Lookup.scala 11:37:@251.4]
  assign _T_210 = _T_74 ? 1'h1 : _T_209; // @[Lookup.scala 11:37:@252.4]
  assign _T_211 = _T_70 ? 1'h1 : _T_210; // @[Lookup.scala 11:37:@253.4]
  assign _T_212 = _T_66 ? 1'h1 : _T_211; // @[Lookup.scala 11:37:@254.4]
  assign _T_213 = _T_62 ? 1'h1 : _T_212; // @[Lookup.scala 11:37:@255.4]
  assign _T_214 = _T_58 ? 1'h1 : _T_213; // @[Lookup.scala 11:37:@256.4]
  assign _T_215 = _T_54 ? 1'h1 : _T_214; // @[Lookup.scala 11:37:@257.4]
  assign _T_216 = _T_50 ? 1'h1 : _T_215; // @[Lookup.scala 11:37:@258.4]
  assign _T_217 = _T_46 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@259.4]
  assign _T_218 = _T_42 ? 1'h1 : _T_217; // @[Lookup.scala 11:37:@260.4]
  assign _T_219 = _T_38 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@261.4]
  assign _T_221 = _T_178 ? 3'h5 : 3'h0; // @[Lookup.scala 11:37:@264.4]
  assign _T_222 = _T_174 ? 3'h5 : _T_221; // @[Lookup.scala 11:37:@265.4]
  assign _T_223 = _T_170 ? 3'h2 : _T_222; // @[Lookup.scala 11:37:@266.4]
  assign _T_224 = _T_166 ? 3'h6 : _T_223; // @[Lookup.scala 11:37:@267.4]
  assign _T_225 = _T_162 ? 3'h4 : _T_224; // @[Lookup.scala 11:37:@268.4]
  assign _T_226 = _T_158 ? 3'h4 : _T_225; // @[Lookup.scala 11:37:@269.4]
  assign _T_227 = _T_154 ? 3'h4 : _T_226; // @[Lookup.scala 11:37:@270.4]
  assign _T_228 = _T_150 ? 3'h4 : _T_227; // @[Lookup.scala 11:37:@271.4]
  assign _T_229 = _T_146 ? 3'h4 : _T_228; // @[Lookup.scala 11:37:@272.4]
  assign _T_230 = _T_142 ? 3'h4 : _T_229; // @[Lookup.scala 11:37:@273.4]
  assign _T_231 = _T_138 ? 3'h3 : _T_230; // @[Lookup.scala 11:37:@274.4]
  assign _T_232 = _T_134 ? 3'h3 : _T_231; // @[Lookup.scala 11:37:@275.4]
  assign _T_233 = _T_130 ? 3'h3 : _T_232; // @[Lookup.scala 11:37:@276.4]
  assign _T_234 = _T_126 ? 3'h2 : _T_233; // @[Lookup.scala 11:37:@277.4]
  assign _T_235 = _T_122 ? 3'h2 : _T_234; // @[Lookup.scala 11:37:@278.4]
  assign _T_236 = _T_118 ? 3'h2 : _T_235; // @[Lookup.scala 11:37:@279.4]
  assign _T_237 = _T_114 ? 3'h2 : _T_236; // @[Lookup.scala 11:37:@280.4]
  assign _T_238 = _T_110 ? 3'h2 : _T_237; // @[Lookup.scala 11:37:@281.4]
  assign _T_239 = _T_106 ? 3'h2 : _T_238; // @[Lookup.scala 11:37:@282.4]
  assign _T_240 = _T_102 ? 3'h2 : _T_239; // @[Lookup.scala 11:37:@283.4]
  assign _T_241 = _T_98 ? 3'h1 : _T_240; // @[Lookup.scala 11:37:@284.4]
  assign _T_242 = _T_94 ? 3'h1 : _T_241; // @[Lookup.scala 11:37:@285.4]
  assign _T_243 = _T_90 ? 3'h2 : _T_242; // @[Lookup.scala 11:37:@286.4]
  assign _T_244 = _T_86 ? 3'h2 : _T_243; // @[Lookup.scala 11:37:@287.4]
  assign _T_245 = _T_82 ? 3'h2 : _T_244; // @[Lookup.scala 11:37:@288.4]
  assign _T_246 = _T_78 ? 3'h1 : _T_245; // @[Lookup.scala 11:37:@289.4]
  assign _T_247 = _T_74 ? 3'h1 : _T_246; // @[Lookup.scala 11:37:@290.4]
  assign _T_248 = _T_70 ? 3'h1 : _T_247; // @[Lookup.scala 11:37:@291.4]
  assign _T_249 = _T_66 ? 3'h2 : _T_248; // @[Lookup.scala 11:37:@292.4]
  assign _T_250 = _T_62 ? 3'h2 : _T_249; // @[Lookup.scala 11:37:@293.4]
  assign _T_251 = _T_58 ? 3'h2 : _T_250; // @[Lookup.scala 11:37:@294.4]
  assign _T_252 = _T_54 ? 3'h2 : _T_251; // @[Lookup.scala 11:37:@295.4]
  assign _T_253 = _T_50 ? 3'h1 : _T_252; // @[Lookup.scala 11:37:@296.4]
  assign _T_254 = _T_46 ? 3'h1 : _T_253; // @[Lookup.scala 11:37:@297.4]
  assign _T_255 = _T_42 ? 3'h1 : _T_254; // @[Lookup.scala 11:37:@298.4]
  assign _T_256 = _T_38 ? 3'h1 : _T_255; // @[Lookup.scala 11:37:@299.4]
  assign _T_269 = _T_134 ? 1'h1 : _T_138; // @[Lookup.scala 11:37:@313.4]
  assign _T_270 = _T_130 ? 1'h1 : _T_269; // @[Lookup.scala 11:37:@314.4]
  assign _T_271 = _T_126 ? 1'h1 : _T_270; // @[Lookup.scala 11:37:@315.4]
  assign _T_272 = _T_122 ? 1'h1 : _T_271; // @[Lookup.scala 11:37:@316.4]
  assign _T_273 = _T_118 ? 1'h1 : _T_272; // @[Lookup.scala 11:37:@317.4]
  assign _T_274 = _T_114 ? 1'h1 : _T_273; // @[Lookup.scala 11:37:@318.4]
  assign _T_275 = _T_110 ? 1'h1 : _T_274; // @[Lookup.scala 11:37:@319.4]
  assign _T_276 = _T_106 ? 1'h1 : _T_275; // @[Lookup.scala 11:37:@320.4]
  assign _T_277 = _T_102 ? 1'h1 : _T_276; // @[Lookup.scala 11:37:@321.4]
  assign _T_278 = _T_98 ? 1'h0 : _T_277; // @[Lookup.scala 11:37:@322.4]
  assign _T_279 = _T_94 ? 1'h0 : _T_278; // @[Lookup.scala 11:37:@323.4]
  assign _T_280 = _T_90 ? 1'h1 : _T_279; // @[Lookup.scala 11:37:@324.4]
  assign _T_281 = _T_86 ? 1'h1 : _T_280; // @[Lookup.scala 11:37:@325.4]
  assign _T_282 = _T_82 ? 1'h1 : _T_281; // @[Lookup.scala 11:37:@326.4]
  assign _T_283 = _T_78 ? 1'h0 : _T_282; // @[Lookup.scala 11:37:@327.4]
  assign _T_284 = _T_74 ? 1'h0 : _T_283; // @[Lookup.scala 11:37:@328.4]
  assign _T_285 = _T_70 ? 1'h0 : _T_284; // @[Lookup.scala 11:37:@329.4]
  assign _T_286 = _T_66 ? 1'h1 : _T_285; // @[Lookup.scala 11:37:@330.4]
  assign _T_287 = _T_62 ? 1'h1 : _T_286; // @[Lookup.scala 11:37:@331.4]
  assign _T_288 = _T_58 ? 1'h1 : _T_287; // @[Lookup.scala 11:37:@332.4]
  assign _T_289 = _T_54 ? 1'h1 : _T_288; // @[Lookup.scala 11:37:@333.4]
  assign _T_290 = _T_50 ? 1'h0 : _T_289; // @[Lookup.scala 11:37:@334.4]
  assign _T_291 = _T_46 ? 1'h0 : _T_290; // @[Lookup.scala 11:37:@335.4]
  assign _T_292 = _T_42 ? 1'h0 : _T_291; // @[Lookup.scala 11:37:@336.4]
  assign _T_293 = _T_38 ? 1'h0 : _T_292; // @[Lookup.scala 11:37:@337.4]
  assign _T_295 = _T_178 ? 5'h0 : 5'h10; // @[Lookup.scala 11:37:@340.4]
  assign _T_296 = _T_174 ? 5'h0 : _T_295; // @[Lookup.scala 11:37:@341.4]
  assign _T_297 = _T_170 ? 5'h0 : _T_296; // @[Lookup.scala 11:37:@342.4]
  assign _T_298 = _T_166 ? 5'h0 : _T_297; // @[Lookup.scala 11:37:@343.4]
  assign _T_299 = _T_162 ? 5'hf : _T_298; // @[Lookup.scala 11:37:@344.4]
  assign _T_300 = _T_158 ? 5'he : _T_299; // @[Lookup.scala 11:37:@345.4]
  assign _T_301 = _T_154 ? 5'hd : _T_300; // @[Lookup.scala 11:37:@346.4]
  assign _T_302 = _T_150 ? 5'hc : _T_301; // @[Lookup.scala 11:37:@347.4]
  assign _T_303 = _T_146 ? 5'hb : _T_302; // @[Lookup.scala 11:37:@348.4]
  assign _T_304 = _T_142 ? 5'ha : _T_303; // @[Lookup.scala 11:37:@349.4]
  assign _T_305 = _T_138 ? 5'h0 : _T_304; // @[Lookup.scala 11:37:@350.4]
  assign _T_306 = _T_134 ? 5'h0 : _T_305; // @[Lookup.scala 11:37:@351.4]
  assign _T_307 = _T_130 ? 5'h0 : _T_306; // @[Lookup.scala 11:37:@352.4]
  assign _T_308 = _T_126 ? 5'h0 : _T_307; // @[Lookup.scala 11:37:@353.4]
  assign _T_309 = _T_122 ? 5'h0 : _T_308; // @[Lookup.scala 11:37:@354.4]
  assign _T_310 = _T_118 ? 5'h0 : _T_309; // @[Lookup.scala 11:37:@355.4]
  assign _T_311 = _T_114 ? 5'h0 : _T_310; // @[Lookup.scala 11:37:@356.4]
  assign _T_312 = _T_110 ? 5'h0 : _T_311; // @[Lookup.scala 11:37:@357.4]
  assign _T_313 = _T_106 ? 5'h9 : _T_312; // @[Lookup.scala 11:37:@358.4]
  assign _T_314 = _T_102 ? 5'h8 : _T_313; // @[Lookup.scala 11:37:@359.4]
  assign _T_315 = _T_98 ? 5'h9 : _T_314; // @[Lookup.scala 11:37:@360.4]
  assign _T_316 = _T_94 ? 5'h8 : _T_315; // @[Lookup.scala 11:37:@361.4]
  assign _T_317 = _T_90 ? 5'h7 : _T_316; // @[Lookup.scala 11:37:@362.4]
  assign _T_318 = _T_86 ? 5'h6 : _T_317; // @[Lookup.scala 11:37:@363.4]
  assign _T_319 = _T_82 ? 5'h5 : _T_318; // @[Lookup.scala 11:37:@364.4]
  assign _T_320 = _T_78 ? 5'h7 : _T_319; // @[Lookup.scala 11:37:@365.4]
  assign _T_321 = _T_74 ? 5'h6 : _T_320; // @[Lookup.scala 11:37:@366.4]
  assign _T_322 = _T_70 ? 5'h5 : _T_321; // @[Lookup.scala 11:37:@367.4]
  assign _T_323 = _T_66 ? 5'h4 : _T_322; // @[Lookup.scala 11:37:@368.4]
  assign _T_324 = _T_62 ? 5'h3 : _T_323; // @[Lookup.scala 11:37:@369.4]
  assign _T_325 = _T_58 ? 5'h2 : _T_324; // @[Lookup.scala 11:37:@370.4]
  assign _T_326 = _T_54 ? 5'h0 : _T_325; // @[Lookup.scala 11:37:@371.4]
  assign _T_327 = _T_50 ? 5'h4 : _T_326; // @[Lookup.scala 11:37:@372.4]
  assign _T_328 = _T_46 ? 5'h3 : _T_327; // @[Lookup.scala 11:37:@373.4]
  assign _T_329 = _T_42 ? 5'h2 : _T_328; // @[Lookup.scala 11:37:@374.4]
  assign _T_330 = _T_38 ? 5'h1 : _T_329; // @[Lookup.scala 11:37:@375.4]
  assign _T_335 = _T_166 ? 1'h1 : _T_170; // @[Lookup.scala 11:37:@381.4]
  assign _T_336 = _T_162 ? 1'h1 : _T_335; // @[Lookup.scala 11:37:@382.4]
  assign _T_337 = _T_158 ? 1'h1 : _T_336; // @[Lookup.scala 11:37:@383.4]
  assign _T_338 = _T_154 ? 1'h1 : _T_337; // @[Lookup.scala 11:37:@384.4]
  assign _T_339 = _T_150 ? 1'h1 : _T_338; // @[Lookup.scala 11:37:@385.4]
  assign _T_340 = _T_146 ? 1'h1 : _T_339; // @[Lookup.scala 11:37:@386.4]
  assign _T_341 = _T_142 ? 1'h1 : _T_340; // @[Lookup.scala 11:37:@387.4]
  assign _T_342 = _T_138 ? 1'h0 : _T_341; // @[Lookup.scala 11:37:@388.4]
  assign _T_343 = _T_134 ? 1'h0 : _T_342; // @[Lookup.scala 11:37:@389.4]
  assign _T_344 = _T_130 ? 1'h0 : _T_343; // @[Lookup.scala 11:37:@390.4]
  assign _T_345 = _T_126 ? 1'h0 : _T_344; // @[Lookup.scala 11:37:@391.4]
  assign _T_346 = _T_122 ? 1'h0 : _T_345; // @[Lookup.scala 11:37:@392.4]
  assign _T_347 = _T_118 ? 1'h0 : _T_346; // @[Lookup.scala 11:37:@393.4]
  assign _T_348 = _T_114 ? 1'h0 : _T_347; // @[Lookup.scala 11:37:@394.4]
  assign _T_349 = _T_110 ? 1'h0 : _T_348; // @[Lookup.scala 11:37:@395.4]
  assign _T_350 = _T_106 ? 1'h0 : _T_349; // @[Lookup.scala 11:37:@396.4]
  assign _T_351 = _T_102 ? 1'h0 : _T_350; // @[Lookup.scala 11:37:@397.4]
  assign _T_352 = _T_98 ? 1'h0 : _T_351; // @[Lookup.scala 11:37:@398.4]
  assign _T_353 = _T_94 ? 1'h0 : _T_352; // @[Lookup.scala 11:37:@399.4]
  assign _T_354 = _T_90 ? 1'h0 : _T_353; // @[Lookup.scala 11:37:@400.4]
  assign _T_355 = _T_86 ? 1'h0 : _T_354; // @[Lookup.scala 11:37:@401.4]
  assign _T_356 = _T_82 ? 1'h0 : _T_355; // @[Lookup.scala 11:37:@402.4]
  assign _T_357 = _T_78 ? 1'h0 : _T_356; // @[Lookup.scala 11:37:@403.4]
  assign _T_358 = _T_74 ? 1'h0 : _T_357; // @[Lookup.scala 11:37:@404.4]
  assign _T_359 = _T_70 ? 1'h0 : _T_358; // @[Lookup.scala 11:37:@405.4]
  assign _T_360 = _T_66 ? 1'h0 : _T_359; // @[Lookup.scala 11:37:@406.4]
  assign _T_361 = _T_62 ? 1'h0 : _T_360; // @[Lookup.scala 11:37:@407.4]
  assign _T_362 = _T_58 ? 1'h0 : _T_361; // @[Lookup.scala 11:37:@408.4]
  assign _T_363 = _T_54 ? 1'h0 : _T_362; // @[Lookup.scala 11:37:@409.4]
  assign _T_364 = _T_50 ? 1'h0 : _T_363; // @[Lookup.scala 11:37:@410.4]
  assign _T_365 = _T_46 ? 1'h0 : _T_364; // @[Lookup.scala 11:37:@411.4]
  assign _T_366 = _T_42 ? 1'h0 : _T_365; // @[Lookup.scala 11:37:@412.4]
  assign _T_367 = _T_38 ? 1'h0 : _T_366; // @[Lookup.scala 11:37:@413.4]
  assign _T_372 = _T_166 ? 1'h0 : _T_170; // @[Lookup.scala 11:37:@419.4]
  assign _T_373 = _T_162 ? 1'h0 : _T_372; // @[Lookup.scala 11:37:@420.4]
  assign _T_374 = _T_158 ? 1'h0 : _T_373; // @[Lookup.scala 11:37:@421.4]
  assign _T_375 = _T_154 ? 1'h0 : _T_374; // @[Lookup.scala 11:37:@422.4]
  assign _T_376 = _T_150 ? 1'h0 : _T_375; // @[Lookup.scala 11:37:@423.4]
  assign _T_377 = _T_146 ? 1'h0 : _T_376; // @[Lookup.scala 11:37:@424.4]
  assign _T_378 = _T_142 ? 1'h0 : _T_377; // @[Lookup.scala 11:37:@425.4]
  assign _T_379 = _T_138 ? 1'h0 : _T_378; // @[Lookup.scala 11:37:@426.4]
  assign _T_380 = _T_134 ? 1'h0 : _T_379; // @[Lookup.scala 11:37:@427.4]
  assign _T_381 = _T_130 ? 1'h0 : _T_380; // @[Lookup.scala 11:37:@428.4]
  assign _T_382 = _T_126 ? 1'h0 : _T_381; // @[Lookup.scala 11:37:@429.4]
  assign _T_383 = _T_122 ? 1'h0 : _T_382; // @[Lookup.scala 11:37:@430.4]
  assign _T_384 = _T_118 ? 1'h0 : _T_383; // @[Lookup.scala 11:37:@431.4]
  assign _T_385 = _T_114 ? 1'h0 : _T_384; // @[Lookup.scala 11:37:@432.4]
  assign _T_386 = _T_110 ? 1'h0 : _T_385; // @[Lookup.scala 11:37:@433.4]
  assign _T_387 = _T_106 ? 1'h0 : _T_386; // @[Lookup.scala 11:37:@434.4]
  assign _T_388 = _T_102 ? 1'h0 : _T_387; // @[Lookup.scala 11:37:@435.4]
  assign _T_389 = _T_98 ? 1'h0 : _T_388; // @[Lookup.scala 11:37:@436.4]
  assign _T_390 = _T_94 ? 1'h0 : _T_389; // @[Lookup.scala 11:37:@437.4]
  assign _T_391 = _T_90 ? 1'h0 : _T_390; // @[Lookup.scala 11:37:@438.4]
  assign _T_392 = _T_86 ? 1'h0 : _T_391; // @[Lookup.scala 11:37:@439.4]
  assign _T_393 = _T_82 ? 1'h0 : _T_392; // @[Lookup.scala 11:37:@440.4]
  assign _T_394 = _T_78 ? 1'h0 : _T_393; // @[Lookup.scala 11:37:@441.4]
  assign _T_395 = _T_74 ? 1'h0 : _T_394; // @[Lookup.scala 11:37:@442.4]
  assign _T_396 = _T_70 ? 1'h0 : _T_395; // @[Lookup.scala 11:37:@443.4]
  assign _T_397 = _T_66 ? 1'h0 : _T_396; // @[Lookup.scala 11:37:@444.4]
  assign _T_398 = _T_62 ? 1'h0 : _T_397; // @[Lookup.scala 11:37:@445.4]
  assign _T_399 = _T_58 ? 1'h0 : _T_398; // @[Lookup.scala 11:37:@446.4]
  assign _T_400 = _T_54 ? 1'h0 : _T_399; // @[Lookup.scala 11:37:@447.4]
  assign _T_401 = _T_50 ? 1'h0 : _T_400; // @[Lookup.scala 11:37:@448.4]
  assign _T_402 = _T_46 ? 1'h0 : _T_401; // @[Lookup.scala 11:37:@449.4]
  assign _T_403 = _T_42 ? 1'h0 : _T_402; // @[Lookup.scala 11:37:@450.4]
  assign _T_404 = _T_38 ? 1'h0 : _T_403; // @[Lookup.scala 11:37:@451.4]
  assign _T_420 = _T_122 ? 1'h1 : _T_126; // @[Lookup.scala 11:37:@468.4]
  assign _T_421 = _T_118 ? 1'h1 : _T_420; // @[Lookup.scala 11:37:@469.4]
  assign _T_422 = _T_114 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@470.4]
  assign _T_423 = _T_110 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@471.4]
  assign _T_424 = _T_106 ? 1'h0 : _T_423; // @[Lookup.scala 11:37:@472.4]
  assign _T_425 = _T_102 ? 1'h0 : _T_424; // @[Lookup.scala 11:37:@473.4]
  assign _T_426 = _T_98 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@474.4]
  assign _T_427 = _T_94 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:@475.4]
  assign _T_428 = _T_90 ? 1'h0 : _T_427; // @[Lookup.scala 11:37:@476.4]
  assign _T_429 = _T_86 ? 1'h0 : _T_428; // @[Lookup.scala 11:37:@477.4]
  assign _T_430 = _T_82 ? 1'h0 : _T_429; // @[Lookup.scala 11:37:@478.4]
  assign _T_431 = _T_78 ? 1'h0 : _T_430; // @[Lookup.scala 11:37:@479.4]
  assign _T_432 = _T_74 ? 1'h0 : _T_431; // @[Lookup.scala 11:37:@480.4]
  assign _T_433 = _T_70 ? 1'h0 : _T_432; // @[Lookup.scala 11:37:@481.4]
  assign _T_434 = _T_66 ? 1'h0 : _T_433; // @[Lookup.scala 11:37:@482.4]
  assign _T_435 = _T_62 ? 1'h0 : _T_434; // @[Lookup.scala 11:37:@483.4]
  assign _T_436 = _T_58 ? 1'h0 : _T_435; // @[Lookup.scala 11:37:@484.4]
  assign _T_437 = _T_54 ? 1'h0 : _T_436; // @[Lookup.scala 11:37:@485.4]
  assign _T_438 = _T_50 ? 1'h0 : _T_437; // @[Lookup.scala 11:37:@486.4]
  assign _T_439 = _T_46 ? 1'h0 : _T_438; // @[Lookup.scala 11:37:@487.4]
  assign _T_440 = _T_42 ? 1'h0 : _T_439; // @[Lookup.scala 11:37:@488.4]
  assign _T_441 = _T_38 ? 1'h0 : _T_440; // @[Lookup.scala 11:37:@489.4]
  assign _T_456 = _T_126 ? 1'h0 : _T_270; // @[Lookup.scala 11:37:@505.4]
  assign _T_457 = _T_122 ? 1'h0 : _T_456; // @[Lookup.scala 11:37:@506.4]
  assign _T_458 = _T_118 ? 1'h0 : _T_457; // @[Lookup.scala 11:37:@507.4]
  assign _T_459 = _T_114 ? 1'h0 : _T_458; // @[Lookup.scala 11:37:@508.4]
  assign _T_460 = _T_110 ? 1'h0 : _T_459; // @[Lookup.scala 11:37:@509.4]
  assign _T_461 = _T_106 ? 1'h0 : _T_460; // @[Lookup.scala 11:37:@510.4]
  assign _T_462 = _T_102 ? 1'h0 : _T_461; // @[Lookup.scala 11:37:@511.4]
  assign _T_463 = _T_98 ? 1'h0 : _T_462; // @[Lookup.scala 11:37:@512.4]
  assign _T_464 = _T_94 ? 1'h0 : _T_463; // @[Lookup.scala 11:37:@513.4]
  assign _T_465 = _T_90 ? 1'h0 : _T_464; // @[Lookup.scala 11:37:@514.4]
  assign _T_466 = _T_86 ? 1'h0 : _T_465; // @[Lookup.scala 11:37:@515.4]
  assign _T_467 = _T_82 ? 1'h0 : _T_466; // @[Lookup.scala 11:37:@516.4]
  assign _T_468 = _T_78 ? 1'h0 : _T_467; // @[Lookup.scala 11:37:@517.4]
  assign _T_469 = _T_74 ? 1'h0 : _T_468; // @[Lookup.scala 11:37:@518.4]
  assign _T_470 = _T_70 ? 1'h0 : _T_469; // @[Lookup.scala 11:37:@519.4]
  assign _T_471 = _T_66 ? 1'h0 : _T_470; // @[Lookup.scala 11:37:@520.4]
  assign _T_472 = _T_62 ? 1'h0 : _T_471; // @[Lookup.scala 11:37:@521.4]
  assign _T_473 = _T_58 ? 1'h0 : _T_472; // @[Lookup.scala 11:37:@522.4]
  assign _T_474 = _T_54 ? 1'h0 : _T_473; // @[Lookup.scala 11:37:@523.4]
  assign _T_475 = _T_50 ? 1'h0 : _T_474; // @[Lookup.scala 11:37:@524.4]
  assign _T_476 = _T_46 ? 1'h0 : _T_475; // @[Lookup.scala 11:37:@525.4]
  assign _T_477 = _T_42 ? 1'h0 : _T_476; // @[Lookup.scala 11:37:@526.4]
  assign _T_478 = _T_38 ? 1'h0 : _T_477; // @[Lookup.scala 11:37:@527.4]
  assign _T_490 = _T_138 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@540.4]
  assign _T_491 = _T_134 ? 2'h1 : _T_490; // @[Lookup.scala 11:37:@541.4]
  assign _T_492 = _T_130 ? 2'h0 : _T_491; // @[Lookup.scala 11:37:@542.4]
  assign _T_493 = _T_126 ? 2'h2 : _T_492; // @[Lookup.scala 11:37:@543.4]
  assign _T_494 = _T_122 ? 2'h1 : _T_493; // @[Lookup.scala 11:37:@544.4]
  assign _T_495 = _T_118 ? 2'h2 : _T_494; // @[Lookup.scala 11:37:@545.4]
  assign _T_496 = _T_114 ? 2'h1 : _T_495; // @[Lookup.scala 11:37:@546.4]
  assign _T_497 = _T_110 ? 2'h0 : _T_496; // @[Lookup.scala 11:37:@547.4]
  assign _T_498 = _T_106 ? 2'h0 : _T_497; // @[Lookup.scala 11:37:@548.4]
  assign _T_499 = _T_102 ? 2'h0 : _T_498; // @[Lookup.scala 11:37:@549.4]
  assign _T_500 = _T_98 ? 2'h0 : _T_499; // @[Lookup.scala 11:37:@550.4]
  assign _T_501 = _T_94 ? 2'h0 : _T_500; // @[Lookup.scala 11:37:@551.4]
  assign _T_502 = _T_90 ? 2'h0 : _T_501; // @[Lookup.scala 11:37:@552.4]
  assign _T_503 = _T_86 ? 2'h0 : _T_502; // @[Lookup.scala 11:37:@553.4]
  assign _T_504 = _T_82 ? 2'h0 : _T_503; // @[Lookup.scala 11:37:@554.4]
  assign _T_505 = _T_78 ? 2'h0 : _T_504; // @[Lookup.scala 11:37:@555.4]
  assign _T_506 = _T_74 ? 2'h0 : _T_505; // @[Lookup.scala 11:37:@556.4]
  assign _T_507 = _T_70 ? 2'h0 : _T_506; // @[Lookup.scala 11:37:@557.4]
  assign _T_508 = _T_66 ? 2'h0 : _T_507; // @[Lookup.scala 11:37:@558.4]
  assign _T_509 = _T_62 ? 2'h0 : _T_508; // @[Lookup.scala 11:37:@559.4]
  assign _T_510 = _T_58 ? 2'h0 : _T_509; // @[Lookup.scala 11:37:@560.4]
  assign _T_511 = _T_54 ? 2'h0 : _T_510; // @[Lookup.scala 11:37:@561.4]
  assign _T_512 = _T_50 ? 2'h0 : _T_511; // @[Lookup.scala 11:37:@562.4]
  assign _T_513 = _T_46 ? 2'h0 : _T_512; // @[Lookup.scala 11:37:@563.4]
  assign _T_514 = _T_42 ? 2'h0 : _T_513; // @[Lookup.scala 11:37:@564.4]
  assign _T_515 = _T_38 ? 2'h0 : _T_514; // @[Lookup.scala 11:37:@565.4]
  assign _T_532 = _T_118 ? 1'h0 : _T_420; // @[Lookup.scala 11:37:@583.4]
  assign _T_533 = _T_114 ? 1'h0 : _T_532; // @[Lookup.scala 11:37:@584.4]
  assign _T_534 = _T_110 ? 1'h0 : _T_533; // @[Lookup.scala 11:37:@585.4]
  assign _T_535 = _T_106 ? 1'h0 : _T_534; // @[Lookup.scala 11:37:@586.4]
  assign _T_536 = _T_102 ? 1'h0 : _T_535; // @[Lookup.scala 11:37:@587.4]
  assign _T_537 = _T_98 ? 1'h0 : _T_536; // @[Lookup.scala 11:37:@588.4]
  assign _T_538 = _T_94 ? 1'h0 : _T_537; // @[Lookup.scala 11:37:@589.4]
  assign _T_539 = _T_90 ? 1'h0 : _T_538; // @[Lookup.scala 11:37:@590.4]
  assign _T_540 = _T_86 ? 1'h0 : _T_539; // @[Lookup.scala 11:37:@591.4]
  assign _T_541 = _T_82 ? 1'h0 : _T_540; // @[Lookup.scala 11:37:@592.4]
  assign _T_542 = _T_78 ? 1'h0 : _T_541; // @[Lookup.scala 11:37:@593.4]
  assign _T_543 = _T_74 ? 1'h0 : _T_542; // @[Lookup.scala 11:37:@594.4]
  assign _T_544 = _T_70 ? 1'h0 : _T_543; // @[Lookup.scala 11:37:@595.4]
  assign _T_545 = _T_66 ? 1'h0 : _T_544; // @[Lookup.scala 11:37:@596.4]
  assign _T_546 = _T_62 ? 1'h0 : _T_545; // @[Lookup.scala 11:37:@597.4]
  assign _T_547 = _T_58 ? 1'h0 : _T_546; // @[Lookup.scala 11:37:@598.4]
  assign _T_548 = _T_54 ? 1'h0 : _T_547; // @[Lookup.scala 11:37:@599.4]
  assign _T_549 = _T_50 ? 1'h0 : _T_548; // @[Lookup.scala 11:37:@600.4]
  assign _T_550 = _T_46 ? 1'h0 : _T_549; // @[Lookup.scala 11:37:@601.4]
  assign _T_551 = _T_42 ? 1'h0 : _T_550; // @[Lookup.scala 11:37:@602.4]
  assign _T_552 = _T_38 ? 1'h0 : _T_551; // @[Lookup.scala 11:37:@603.4]
  assign _T_554 = _T_178 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@606.4]
  assign _T_555 = _T_174 ? 3'h3 : _T_554; // @[Lookup.scala 11:37:@607.4]
  assign _T_556 = _T_170 ? 3'h2 : _T_555; // @[Lookup.scala 11:37:@608.4]
  assign _T_557 = _T_166 ? 3'h2 : _T_556; // @[Lookup.scala 11:37:@609.4]
  assign _T_558 = _T_162 ? 3'h0 : _T_557; // @[Lookup.scala 11:37:@610.4]
  assign _T_559 = _T_158 ? 3'h0 : _T_558; // @[Lookup.scala 11:37:@611.4]
  assign _T_560 = _T_154 ? 3'h0 : _T_559; // @[Lookup.scala 11:37:@612.4]
  assign _T_561 = _T_150 ? 3'h0 : _T_560; // @[Lookup.scala 11:37:@613.4]
  assign _T_562 = _T_146 ? 3'h0 : _T_561; // @[Lookup.scala 11:37:@614.4]
  assign _T_563 = _T_142 ? 3'h0 : _T_562; // @[Lookup.scala 11:37:@615.4]
  assign _T_564 = _T_138 ? 3'h0 : _T_563; // @[Lookup.scala 11:37:@616.4]
  assign _T_565 = _T_134 ? 3'h0 : _T_564; // @[Lookup.scala 11:37:@617.4]
  assign _T_566 = _T_130 ? 3'h0 : _T_565; // @[Lookup.scala 11:37:@618.4]
  assign _T_567 = _T_126 ? 3'h1 : _T_566; // @[Lookup.scala 11:37:@619.4]
  assign _T_568 = _T_122 ? 3'h1 : _T_567; // @[Lookup.scala 11:37:@620.4]
  assign _T_569 = _T_118 ? 3'h1 : _T_568; // @[Lookup.scala 11:37:@621.4]
  assign _T_570 = _T_114 ? 3'h1 : _T_569; // @[Lookup.scala 11:37:@622.4]
  assign _T_571 = _T_110 ? 3'h1 : _T_570; // @[Lookup.scala 11:37:@623.4]
  assign _T_572 = _T_106 ? 3'h0 : _T_571; // @[Lookup.scala 11:37:@624.4]
  assign _T_573 = _T_102 ? 3'h0 : _T_572; // @[Lookup.scala 11:37:@625.4]
  assign _T_574 = _T_98 ? 3'h0 : _T_573; // @[Lookup.scala 11:37:@626.4]
  assign _T_575 = _T_94 ? 3'h0 : _T_574; // @[Lookup.scala 11:37:@627.4]
  assign _T_576 = _T_90 ? 3'h0 : _T_575; // @[Lookup.scala 11:37:@628.4]
  assign _T_577 = _T_86 ? 3'h0 : _T_576; // @[Lookup.scala 11:37:@629.4]
  assign _T_578 = _T_82 ? 3'h0 : _T_577; // @[Lookup.scala 11:37:@630.4]
  assign _T_579 = _T_78 ? 3'h0 : _T_578; // @[Lookup.scala 11:37:@631.4]
  assign _T_580 = _T_74 ? 3'h0 : _T_579; // @[Lookup.scala 11:37:@632.4]
  assign _T_581 = _T_70 ? 3'h0 : _T_580; // @[Lookup.scala 11:37:@633.4]
  assign _T_582 = _T_66 ? 3'h0 : _T_581; // @[Lookup.scala 11:37:@634.4]
  assign _T_583 = _T_62 ? 3'h0 : _T_582; // @[Lookup.scala 11:37:@635.4]
  assign _T_584 = _T_58 ? 3'h0 : _T_583; // @[Lookup.scala 11:37:@636.4]
  assign _T_585 = _T_54 ? 3'h0 : _T_584; // @[Lookup.scala 11:37:@637.4]
  assign _T_586 = _T_50 ? 3'h0 : _T_585; // @[Lookup.scala 11:37:@638.4]
  assign _T_587 = _T_46 ? 3'h0 : _T_586; // @[Lookup.scala 11:37:@639.4]
  assign _T_588 = _T_42 ? 3'h0 : _T_587; // @[Lookup.scala 11:37:@640.4]
  assign _T_589 = _T_38 ? 3'h0 : _T_588; // @[Lookup.scala 11:37:@641.4]
  assign _T_595 = _T_162 ? 1'h0 : _T_335; // @[Lookup.scala 11:37:@648.4]
  assign _T_596 = _T_158 ? 1'h0 : _T_595; // @[Lookup.scala 11:37:@649.4]
  assign _T_597 = _T_154 ? 1'h0 : _T_596; // @[Lookup.scala 11:37:@650.4]
  assign _T_598 = _T_150 ? 1'h0 : _T_597; // @[Lookup.scala 11:37:@651.4]
  assign _T_599 = _T_146 ? 1'h0 : _T_598; // @[Lookup.scala 11:37:@652.4]
  assign _T_600 = _T_142 ? 1'h0 : _T_599; // @[Lookup.scala 11:37:@653.4]
  assign _T_601 = _T_138 ? 1'h0 : _T_600; // @[Lookup.scala 11:37:@654.4]
  assign _T_602 = _T_134 ? 1'h0 : _T_601; // @[Lookup.scala 11:37:@655.4]
  assign _T_603 = _T_130 ? 1'h0 : _T_602; // @[Lookup.scala 11:37:@656.4]
  assign _T_604 = _T_126 ? 1'h0 : _T_603; // @[Lookup.scala 11:37:@657.4]
  assign _T_605 = _T_122 ? 1'h0 : _T_604; // @[Lookup.scala 11:37:@658.4]
  assign _T_606 = _T_118 ? 1'h0 : _T_605; // @[Lookup.scala 11:37:@659.4]
  assign _T_607 = _T_114 ? 1'h0 : _T_606; // @[Lookup.scala 11:37:@660.4]
  assign _T_608 = _T_110 ? 1'h0 : _T_607; // @[Lookup.scala 11:37:@661.4]
  assign _T_609 = _T_106 ? 1'h0 : _T_608; // @[Lookup.scala 11:37:@662.4]
  assign _T_610 = _T_102 ? 1'h0 : _T_609; // @[Lookup.scala 11:37:@663.4]
  assign _T_611 = _T_98 ? 1'h0 : _T_610; // @[Lookup.scala 11:37:@664.4]
  assign _T_612 = _T_94 ? 1'h0 : _T_611; // @[Lookup.scala 11:37:@665.4]
  assign _T_613 = _T_90 ? 1'h0 : _T_612; // @[Lookup.scala 11:37:@666.4]
  assign _T_614 = _T_86 ? 1'h0 : _T_613; // @[Lookup.scala 11:37:@667.4]
  assign _T_615 = _T_82 ? 1'h0 : _T_614; // @[Lookup.scala 11:37:@668.4]
  assign _T_616 = _T_78 ? 1'h0 : _T_615; // @[Lookup.scala 11:37:@669.4]
  assign _T_617 = _T_74 ? 1'h0 : _T_616; // @[Lookup.scala 11:37:@670.4]
  assign _T_618 = _T_70 ? 1'h0 : _T_617; // @[Lookup.scala 11:37:@671.4]
  assign _T_619 = _T_66 ? 1'h0 : _T_618; // @[Lookup.scala 11:37:@672.4]
  assign _T_620 = _T_62 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@673.4]
  assign _T_621 = _T_58 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@674.4]
  assign _T_622 = _T_54 ? 1'h0 : _T_621; // @[Lookup.scala 11:37:@675.4]
  assign _T_623 = _T_50 ? 1'h0 : _T_622; // @[Lookup.scala 11:37:@676.4]
  assign _T_624 = _T_46 ? 1'h0 : _T_623; // @[Lookup.scala 11:37:@677.4]
  assign _T_625 = _T_42 ? 1'h0 : _T_624; // @[Lookup.scala 11:37:@678.4]
  assign _T_626 = _T_38 ? 1'h0 : _T_625; // @[Lookup.scala 11:37:@679.4]
  assign io_Reg_Write = _T_34 ? 1'h1 : _T_219; // @[Control.scala 174:17:@691.4]
  assign io_Imm_Sel = _T_34 ? 3'h1 : _T_256; // @[Control.scala 158:17:@681.4]
  assign io_ALU_Src = _T_34 ? 1'h0 : _T_293; // @[Control.scala 161:17:@682.4]
  assign io_ALUOp = _T_34 ? 5'h0 : _T_330; // @[Control.scala 162:17:@683.4]
  assign io_Branch = _T_34 ? 1'h0 : _T_367; // @[Control.scala 163:17:@684.4]
  assign io_Branch_Src = _T_34 ? 1'h0 : _T_404; // @[Control.scala 164:17:@685.4]
  assign io_Mem_Read = _T_34 ? 1'h0 : _T_441; // @[Control.scala 168:17:@687.4]
  assign io_Mem_Write = _T_34 ? 1'h0 : _T_478; // @[Control.scala 169:17:@688.4]
  assign io_Data_Size = _T_34 ? 2'h0 : _T_515; // @[Control.scala 170:17:@689.4]
  assign io_Load_Type = _T_34 ? 1'h0 : _T_552; // @[Control.scala 171:17:@690.4]
  assign io_Mem_to_Reg = _T_34 ? 3'h0 : _T_589; // @[Control.scala 175:17:@692.4]
  assign io_Jump_Type = _T_34 ? 1'h0 : _T_626; // @[Control.scala 165:17:@686.4]
endmodule
module ID_EX_Register( // @[:@694.2]
  input         clock, // @[:@695.4]
  input         reset, // @[:@696.4]
  input  [31:0] io_id_pc, // @[:@697.4]
  input  [31:0] io_id_pc_4, // @[:@697.4]
  input  [31:0] io_id_rs1_out, // @[:@697.4]
  input  [31:0] io_id_rs2_out, // @[:@697.4]
  input  [31:0] io_id_imm, // @[:@697.4]
  input  [31:0] io_id_inst, // @[:@697.4]
  input  [4:0]  io_id_rs1, // @[:@697.4]
  input  [4:0]  io_id_rs2, // @[:@697.4]
  input         io_ALU_Src, // @[:@697.4]
  input  [4:0]  io_ALUOp, // @[:@697.4]
  input         io_Branch, // @[:@697.4]
  input         io_Branch_Src, // @[:@697.4]
  input         io_Jump_Type, // @[:@697.4]
  input         io_Mem_Read, // @[:@697.4]
  input         io_Mem_Write, // @[:@697.4]
  input  [1:0]  io_Data_Size, // @[:@697.4]
  input         io_Load_Type, // @[:@697.4]
  input         io_Reg_Write, // @[:@697.4]
  input  [2:0]  io_Mem_to_Reg, // @[:@697.4]
  output        io_ex_ALU_Src, // @[:@697.4]
  output [4:0]  io_ex_ALUOp, // @[:@697.4]
  output        io_ex_Branch, // @[:@697.4]
  output        io_ex_Branch_Src, // @[:@697.4]
  output        io_ex_Jump_Type, // @[:@697.4]
  output        io_ex_Mem_Read, // @[:@697.4]
  output        io_ex_Mem_Write, // @[:@697.4]
  output [1:0]  io_ex_Data_Size, // @[:@697.4]
  output        io_ex_Load_Type, // @[:@697.4]
  output        io_ex_Reg_Write, // @[:@697.4]
  output [2:0]  io_ex_Mem_to_Reg, // @[:@697.4]
  output [31:0] io_ex_pc, // @[:@697.4]
  output [31:0] io_ex_pc_4, // @[:@697.4]
  output [31:0] io_ex_rs1_out, // @[:@697.4]
  output [31:0] io_ex_rs2_out, // @[:@697.4]
  output [4:0]  io_ex_rd, // @[:@697.4]
  output [31:0] io_ex_imm, // @[:@697.4]
  output [4:0]  io_ex_rs1, // @[:@697.4]
  output [4:0]  io_ex_rs2 // @[:@697.4]
);
  reg [31:0] pc; // @[ID_EX_Register.scala 70:28:@699.4]
  reg [31:0] _RAND_0;
  reg [31:0] pc_4; // @[ID_EX_Register.scala 71:28:@700.4]
  reg [31:0] _RAND_1;
  reg [31:0] rs1_out; // @[ID_EX_Register.scala 72:28:@701.4]
  reg [31:0] _RAND_2;
  reg [31:0] rs2_out; // @[ID_EX_Register.scala 73:28:@702.4]
  reg [31:0] _RAND_3;
  reg [31:0] imm; // @[ID_EX_Register.scala 74:28:@703.4]
  reg [31:0] _RAND_4;
  reg [31:0] inst; // @[ID_EX_Register.scala 75:28:@704.4]
  reg [31:0] _RAND_5;
  reg [31:0] rs1; // @[ID_EX_Register.scala 76:28:@705.4]
  reg [31:0] _RAND_6;
  reg [31:0] rs2; // @[ID_EX_Register.scala 77:28:@706.4]
  reg [31:0] _RAND_7;
  reg  alu_src; // @[ID_EX_Register.scala 78:28:@707.4]
  reg [31:0] _RAND_8;
  reg [4:0] aluop; // @[ID_EX_Register.scala 79:28:@708.4]
  reg [31:0] _RAND_9;
  reg  branch; // @[ID_EX_Register.scala 80:28:@709.4]
  reg [31:0] _RAND_10;
  reg  branch_src; // @[ID_EX_Register.scala 81:28:@710.4]
  reg [31:0] _RAND_11;
  reg  jump_type; // @[ID_EX_Register.scala 82:28:@711.4]
  reg [31:0] _RAND_12;
  reg  mem_read; // @[ID_EX_Register.scala 83:28:@712.4]
  reg [31:0] _RAND_13;
  reg  mem_write; // @[ID_EX_Register.scala 84:28:@713.4]
  reg [31:0] _RAND_14;
  reg [1:0] data_size; // @[ID_EX_Register.scala 85:28:@714.4]
  reg [31:0] _RAND_15;
  reg  load_type; // @[ID_EX_Register.scala 86:28:@715.4]
  reg [31:0] _RAND_16;
  reg  reg_write; // @[ID_EX_Register.scala 87:28:@716.4]
  reg [31:0] _RAND_17;
  reg [2:0] mem_to_reg; // @[ID_EX_Register.scala 88:28:@717.4]
  reg [31:0] _RAND_18;
  assign io_ex_ALU_Src = alu_src; // @[ID_EX_Register.scala 112:21:@737.4]
  assign io_ex_ALUOp = aluop; // @[ID_EX_Register.scala 113:21:@738.4]
  assign io_ex_Branch = branch; // @[ID_EX_Register.scala 114:21:@739.4]
  assign io_ex_Branch_Src = branch_src; // @[ID_EX_Register.scala 115:21:@740.4]
  assign io_ex_Jump_Type = jump_type; // @[ID_EX_Register.scala 116:21:@741.4]
  assign io_ex_Mem_Read = mem_read; // @[ID_EX_Register.scala 117:21:@742.4]
  assign io_ex_Mem_Write = mem_write; // @[ID_EX_Register.scala 118:21:@743.4]
  assign io_ex_Data_Size = data_size; // @[ID_EX_Register.scala 121:21:@746.4]
  assign io_ex_Load_Type = load_type; // @[ID_EX_Register.scala 122:21:@747.4]
  assign io_ex_Reg_Write = reg_write; // @[ID_EX_Register.scala 119:21:@744.4]
  assign io_ex_Mem_to_Reg = mem_to_reg; // @[ID_EX_Register.scala 120:21:@745.4]
  assign io_ex_pc = pc; // @[ID_EX_Register.scala 123:21:@748.4]
  assign io_ex_pc_4 = pc_4; // @[ID_EX_Register.scala 124:21:@749.4]
  assign io_ex_rs1_out = rs1_out; // @[ID_EX_Register.scala 125:21:@750.4]
  assign io_ex_rs2_out = rs2_out; // @[ID_EX_Register.scala 126:21:@751.4]
  assign io_ex_rd = inst[11:7]; // @[ID_EX_Register.scala 131:21:@757.4]
  assign io_ex_imm = imm; // @[ID_EX_Register.scala 129:21:@754.4]
  assign io_ex_rs1 = rs1[4:0]; // @[ID_EX_Register.scala 127:21:@752.4]
  assign io_ex_rs2 = rs2[4:0]; // @[ID_EX_Register.scala 128:21:@753.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc_4 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rs1_out = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rs2_out = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imm = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  inst = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rs1 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rs2 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  alu_src = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  aluop = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  branch = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  branch_src = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  jump_type = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_read = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_write = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  data_size = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  load_type = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_write = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_to_reg = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h0;
    end else begin
      pc <= io_id_pc;
    end
    if (reset) begin
      pc_4 <= 32'h0;
    end else begin
      pc_4 <= io_id_pc_4;
    end
    if (reset) begin
      rs1_out <= 32'h0;
    end else begin
      rs1_out <= io_id_rs1_out;
    end
    if (reset) begin
      rs2_out <= 32'h0;
    end else begin
      rs2_out <= io_id_rs2_out;
    end
    if (reset) begin
      imm <= 32'h0;
    end else begin
      imm <= io_id_imm;
    end
    if (reset) begin
      inst <= 32'h0;
    end else begin
      inst <= io_id_inst;
    end
    if (reset) begin
      rs1 <= 32'h0;
    end else begin
      rs1 <= {{27'd0}, io_id_rs1};
    end
    if (reset) begin
      rs2 <= 32'h0;
    end else begin
      rs2 <= {{27'd0}, io_id_rs2};
    end
    if (reset) begin
      alu_src <= 1'h0;
    end else begin
      alu_src <= io_ALU_Src;
    end
    if (reset) begin
      aluop <= 5'h0;
    end else begin
      aluop <= io_ALUOp;
    end
    if (reset) begin
      branch <= 1'h0;
    end else begin
      branch <= io_Branch;
    end
    if (reset) begin
      branch_src <= 1'h0;
    end else begin
      branch_src <= io_Branch_Src;
    end
    if (reset) begin
      jump_type <= 1'h0;
    end else begin
      jump_type <= io_Jump_Type;
    end
    if (reset) begin
      mem_read <= 1'h0;
    end else begin
      mem_read <= io_Mem_Read;
    end
    if (reset) begin
      mem_write <= 1'h0;
    end else begin
      mem_write <= io_Mem_Write;
    end
    if (reset) begin
      data_size <= 2'h0;
    end else begin
      data_size <= io_Data_Size;
    end
    if (reset) begin
      load_type <= 1'h0;
    end else begin
      load_type <= io_Load_Type;
    end
    if (reset) begin
      reg_write <= 1'h0;
    end else begin
      reg_write <= io_Reg_Write;
    end
    if (reset) begin
      mem_to_reg <= 3'h0;
    end else begin
      mem_to_reg <= io_Mem_to_Reg;
    end
  end
endmodule
module ALU( // @[:@759.2]
  input  [31:0] io_Src_A, // @[:@762.4]
  input  [31:0] io_Src_B, // @[:@762.4]
  input  [4:0]  io_ALUOp, // @[:@762.4]
  output [31:0] io_Sum, // @[:@762.4]
  output        io_Conflag // @[:@762.4]
);
  wire [5:0] shamt; // @[ALU.scala 52:23:@764.4]
  wire [32:0] _T_15; // @[ALU.scala 54:28:@765.4]
  wire [31:0] _T_16; // @[ALU.scala 54:28:@766.4]
  wire [32:0] _T_17; // @[ALU.scala 55:28:@767.4]
  wire [32:0] _T_18; // @[ALU.scala 55:28:@768.4]
  wire [31:0] _T_19; // @[ALU.scala 55:28:@769.4]
  wire [31:0] _T_20; // @[ALU.scala 56:28:@770.4]
  wire [31:0] _T_21; // @[ALU.scala 57:28:@771.4]
  wire [31:0] _GEN_0; // @[ALU.scala 58:28:@772.4]
  wire [31:0] _T_22; // @[ALU.scala 58:28:@772.4]
  wire [94:0] _GEN_1; // @[ALU.scala 59:28:@773.4]
  wire [94:0] _T_23; // @[ALU.scala 59:28:@773.4]
  wire [31:0] _T_24; // @[ALU.scala 60:28:@774.4]
  wire [31:0] _T_25; // @[ALU.scala 61:34:@775.4]
  wire [31:0] _T_26; // @[ALU.scala 61:37:@776.4]
  wire [31:0] _T_27; // @[ALU.scala 61:53:@777.4]
  wire [31:0] _T_29; // @[ALU.scala 62:54:@779.4]
  wire  _T_30; // @[ALU.scala 62:37:@780.4]
  wire  _T_31; // @[ALU.scala 63:28:@781.4]
  wire  _T_32; // @[Mux.scala 46:19:@782.4]
  wire [31:0] _T_33; // @[Mux.scala 46:16:@783.4]
  wire  _T_34; // @[Mux.scala 46:19:@784.4]
  wire [31:0] _T_35; // @[Mux.scala 46:16:@785.4]
  wire  _T_36; // @[Mux.scala 46:19:@786.4]
  wire [31:0] _T_37; // @[Mux.scala 46:16:@787.4]
  wire  _T_38; // @[Mux.scala 46:19:@788.4]
  wire [31:0] _T_39; // @[Mux.scala 46:16:@789.4]
  wire  _T_40; // @[Mux.scala 46:19:@790.4]
  wire [94:0] _T_41; // @[Mux.scala 46:16:@791.4]
  wire  _T_42; // @[Mux.scala 46:19:@792.4]
  wire [94:0] _T_43; // @[Mux.scala 46:16:@793.4]
  wire  _T_44; // @[Mux.scala 46:19:@794.4]
  wire [94:0] _T_45; // @[Mux.scala 46:16:@795.4]
  wire  _T_46; // @[Mux.scala 46:19:@796.4]
  wire [94:0] _T_47; // @[Mux.scala 46:16:@797.4]
  wire  _T_48; // @[Mux.scala 46:19:@798.4]
  wire [94:0] _T_49; // @[Mux.scala 46:16:@799.4]
  wire  _T_50; // @[Mux.scala 46:19:@800.4]
  wire [94:0] _T_51; // @[Mux.scala 46:16:@801.4]
  wire  _T_55; // @[ALU.scala 67:37:@805.4]
  wire  _T_58; // @[ALU.scala 68:37:@808.4]
  wire  _T_64; // @[ALU.scala 70:37:@814.4]
  wire  _T_66; // @[ALU.scala 72:28:@816.4]
  wire  _T_67; // @[Mux.scala 46:19:@817.4]
  wire  _T_68; // @[Mux.scala 46:16:@818.4]
  wire  _T_69; // @[Mux.scala 46:19:@819.4]
  wire  _T_70; // @[Mux.scala 46:16:@820.4]
  wire  _T_71; // @[Mux.scala 46:19:@821.4]
  wire  _T_72; // @[Mux.scala 46:16:@822.4]
  wire  _T_73; // @[Mux.scala 46:19:@823.4]
  wire  _T_74; // @[Mux.scala 46:16:@824.4]
  wire  _T_75; // @[Mux.scala 46:19:@825.4]
  wire  _T_76; // @[Mux.scala 46:16:@826.4]
  wire  _T_77; // @[Mux.scala 46:19:@827.4]
  assign shamt = io_Src_B[5:0]; // @[ALU.scala 52:23:@764.4]
  assign _T_15 = io_Src_A + io_Src_B; // @[ALU.scala 54:28:@765.4]
  assign _T_16 = io_Src_A + io_Src_B; // @[ALU.scala 54:28:@766.4]
  assign _T_17 = io_Src_A - io_Src_B; // @[ALU.scala 55:28:@767.4]
  assign _T_18 = $unsigned(_T_17); // @[ALU.scala 55:28:@768.4]
  assign _T_19 = _T_18[31:0]; // @[ALU.scala 55:28:@769.4]
  assign _T_20 = io_Src_A & io_Src_B; // @[ALU.scala 56:28:@770.4]
  assign _T_21 = io_Src_A | io_Src_B; // @[ALU.scala 57:28:@771.4]
  assign _GEN_0 = {{26'd0}, shamt}; // @[ALU.scala 58:28:@772.4]
  assign _T_22 = io_Src_A ^ _GEN_0; // @[ALU.scala 58:28:@772.4]
  assign _GEN_1 = {{63'd0}, io_Src_A}; // @[ALU.scala 59:28:@773.4]
  assign _T_23 = _GEN_1 << shamt; // @[ALU.scala 59:28:@773.4]
  assign _T_24 = io_Src_A >> shamt; // @[ALU.scala 60:28:@774.4]
  assign _T_25 = $signed(io_Src_A); // @[ALU.scala 61:34:@775.4]
  assign _T_26 = $signed(_T_25) >>> shamt; // @[ALU.scala 61:37:@776.4]
  assign _T_27 = $unsigned(_T_26); // @[ALU.scala 61:53:@777.4]
  assign _T_29 = $signed(io_Src_B); // @[ALU.scala 62:54:@779.4]
  assign _T_30 = $signed(_T_25) < $signed(_T_29); // @[ALU.scala 62:37:@780.4]
  assign _T_31 = io_Src_A < io_Src_B; // @[ALU.scala 63:28:@781.4]
  assign _T_32 = 5'h9 == io_ALUOp; // @[Mux.scala 46:19:@782.4]
  assign _T_33 = _T_32 ? {{31'd0}, _T_31} : io_Src_B; // @[Mux.scala 46:16:@783.4]
  assign _T_34 = 5'h8 == io_ALUOp; // @[Mux.scala 46:19:@784.4]
  assign _T_35 = _T_34 ? {{31'd0}, _T_30} : _T_33; // @[Mux.scala 46:16:@785.4]
  assign _T_36 = 5'h7 == io_ALUOp; // @[Mux.scala 46:19:@786.4]
  assign _T_37 = _T_36 ? _T_27 : _T_35; // @[Mux.scala 46:16:@787.4]
  assign _T_38 = 5'h6 == io_ALUOp; // @[Mux.scala 46:19:@788.4]
  assign _T_39 = _T_38 ? _T_24 : _T_37; // @[Mux.scala 46:16:@789.4]
  assign _T_40 = 5'h5 == io_ALUOp; // @[Mux.scala 46:19:@790.4]
  assign _T_41 = _T_40 ? _T_23 : {{63'd0}, _T_39}; // @[Mux.scala 46:16:@791.4]
  assign _T_42 = 5'h4 == io_ALUOp; // @[Mux.scala 46:19:@792.4]
  assign _T_43 = _T_42 ? {{63'd0}, _T_22} : _T_41; // @[Mux.scala 46:16:@793.4]
  assign _T_44 = 5'h3 == io_ALUOp; // @[Mux.scala 46:19:@794.4]
  assign _T_45 = _T_44 ? {{63'd0}, _T_21} : _T_43; // @[Mux.scala 46:16:@795.4]
  assign _T_46 = 5'h2 == io_ALUOp; // @[Mux.scala 46:19:@796.4]
  assign _T_47 = _T_46 ? {{63'd0}, _T_20} : _T_45; // @[Mux.scala 46:16:@797.4]
  assign _T_48 = 5'h1 == io_ALUOp; // @[Mux.scala 46:19:@798.4]
  assign _T_49 = _T_48 ? {{63'd0}, _T_19} : _T_47; // @[Mux.scala 46:16:@799.4]
  assign _T_50 = 5'h0 == io_ALUOp; // @[Mux.scala 46:19:@800.4]
  assign _T_51 = _T_50 ? {{63'd0}, _T_16} : _T_49; // @[Mux.scala 46:16:@801.4]
  assign _T_55 = $signed(_T_25) == $signed(_T_29); // @[ALU.scala 67:37:@805.4]
  assign _T_58 = $signed(_T_25) != $signed(_T_29); // @[ALU.scala 68:37:@808.4]
  assign _T_64 = $signed(_T_25) >= $signed(_T_29); // @[ALU.scala 70:37:@814.4]
  assign _T_66 = io_Src_A >= io_Src_B; // @[ALU.scala 72:28:@816.4]
  assign _T_67 = 5'hf == io_ALUOp; // @[Mux.scala 46:19:@817.4]
  assign _T_68 = _T_67 ? _T_66 : 1'h0; // @[Mux.scala 46:16:@818.4]
  assign _T_69 = 5'he == io_ALUOp; // @[Mux.scala 46:19:@819.4]
  assign _T_70 = _T_69 ? _T_31 : _T_68; // @[Mux.scala 46:16:@820.4]
  assign _T_71 = 5'hd == io_ALUOp; // @[Mux.scala 46:19:@821.4]
  assign _T_72 = _T_71 ? _T_64 : _T_70; // @[Mux.scala 46:16:@822.4]
  assign _T_73 = 5'hc == io_ALUOp; // @[Mux.scala 46:19:@823.4]
  assign _T_74 = _T_73 ? _T_30 : _T_72; // @[Mux.scala 46:16:@824.4]
  assign _T_75 = 5'hb == io_ALUOp; // @[Mux.scala 46:19:@825.4]
  assign _T_76 = _T_75 ? _T_58 : _T_74; // @[Mux.scala 46:16:@826.4]
  assign _T_77 = 5'ha == io_ALUOp; // @[Mux.scala 46:19:@827.4]
  assign io_Sum = _T_51[31:0]; // @[ALU.scala 53:10:@802.4]
  assign io_Conflag = _T_77 ? _T_55 : _T_76; // @[ALU.scala 66:14:@829.4]
endmodule
module Datapath( // @[:@831.2]
  input  [31:0] io_if_datapathio_if_pc, // @[:@834.4]
  output [31:0] io_if_datapathio_if_new_pc, // @[:@834.4]
  output [31:0] io_if_datapathio_if_pc_4, // @[:@834.4]
  input  [31:0] io_ex_datapathio_ex_rs1_out, // @[:@834.4]
  input  [31:0] io_ex_datapathio_ex_rs2_out, // @[:@834.4]
  input  [31:0] io_ex_datapathio_ex_imm, // @[:@834.4]
  input  [31:0] io_ex_datapathio_ex_pc, // @[:@834.4]
  input         io_ex_datapathio_ex_ALU_Src, // @[:@834.4]
  input         io_ex_datapathio_ex_Branch, // @[:@834.4]
  input         io_ex_datapathio_ex_alu_conflag, // @[:@834.4]
  input         io_ex_datapathio_ex_Branch_Src, // @[:@834.4]
  input         io_ex_datapathio_ex_Jump_Type, // @[:@834.4]
  input  [31:0] io_ex_datapathio_mem_alu_sum, // @[:@834.4]
  input  [1:0]  io_ex_datapathio_Forward_A, // @[:@834.4]
  input  [1:0]  io_ex_datapathio_Forward_B, // @[:@834.4]
  output [31:0] io_ex_datapathio_alu_b_src, // @[:@834.4]
  output [31:0] io_ex_datapathio_ex_aui_pc, // @[:@834.4]
  output [31:0] io_ex_datapathio_forward_rs2_out, // @[:@834.4]
  output [31:0] io_ex_datapathio_alu_a_src, // @[:@834.4]
  input  [31:0] io_wb_datapathio_wb_alu_sum, // @[:@834.4]
  input  [31:0] io_wb_datapathio_wb_dataout, // @[:@834.4]
  input  [31:0] io_wb_datapathio_wb_pc_4, // @[:@834.4]
  input  [31:0] io_wb_datapathio_wb_imm, // @[:@834.4]
  input  [31:0] io_wb_datapathio_wb_aui_pc, // @[:@834.4]
  input  [2:0]  io_wb_datapathio_wb_Mem_to_Reg, // @[:@834.4]
  output [31:0] io_wb_datapathio_wb_reg_writedata // @[:@834.4]
);
  wire [32:0] _T_58; // @[Datapath.scala 66:37:@836.4]
  wire [31:0] PC_4; // @[Datapath.scala 66:37:@837.4]
  wire [31:0] _T_60; // @[Datapath.scala 70:27:@840.4]
  wire [32:0] _T_61; // @[Datapath.scala 70:121:@841.4]
  wire [31:0] ex_branch_addr; // @[Datapath.scala 70:121:@842.4]
  wire  _T_64; // @[Datapath.scala 75:19:@845.4]
  wire  PC_Src; // @[Datapath.scala 75:98:@846.4]
  wire  _T_73; // @[Mux.scala 46:19:@850.4]
  wire [31:0] _T_74; // @[Mux.scala 46:16:@851.4]
  wire  _T_75; // @[Mux.scala 46:19:@852.4]
  wire [31:0] _T_76; // @[Mux.scala 46:16:@853.4]
  wire  _T_77; // @[Mux.scala 46:19:@854.4]
  wire  _T_79; // @[Mux.scala 46:19:@857.4]
  wire [31:0] _T_80; // @[Mux.scala 46:16:@858.4]
  wire  _T_81; // @[Mux.scala 46:19:@859.4]
  wire [31:0] _T_82; // @[Mux.scala 46:16:@860.4]
  wire  _T_83; // @[Mux.scala 46:19:@861.4]
  wire [31:0] operand_b; // @[Mux.scala 46:16:@862.4]
  wire  _T_86; // @[Mux.scala 46:19:@867.4]
  wire [31:0] _T_87; // @[Mux.scala 46:16:@868.4]
  wire  _T_88; // @[Mux.scala 46:19:@869.4]
  wire [31:0] _T_89; // @[Mux.scala 46:16:@870.4]
  wire  _T_90; // @[Mux.scala 46:19:@871.4]
  wire [31:0] _T_91; // @[Mux.scala 46:16:@872.4]
  wire  _T_92; // @[Mux.scala 46:19:@873.4]
  wire [31:0] _T_93; // @[Mux.scala 46:16:@874.4]
  wire  _T_94; // @[Mux.scala 46:19:@875.4]
  assign _T_58 = io_if_datapathio_if_pc + 32'h4; // @[Datapath.scala 66:37:@836.4]
  assign PC_4 = io_if_datapathio_if_pc + 32'h4; // @[Datapath.scala 66:37:@837.4]
  assign _T_60 = io_ex_datapathio_ex_Branch_Src ? io_ex_datapathio_alu_a_src : io_ex_datapathio_ex_pc; // @[Datapath.scala 70:27:@840.4]
  assign _T_61 = _T_60 + io_ex_datapathio_ex_imm; // @[Datapath.scala 70:121:@841.4]
  assign ex_branch_addr = _T_60 + io_ex_datapathio_ex_imm; // @[Datapath.scala 70:121:@842.4]
  assign _T_64 = io_ex_datapathio_ex_Jump_Type ? 1'h1 : io_ex_datapathio_ex_alu_conflag; // @[Datapath.scala 75:19:@845.4]
  assign PC_Src = _T_64 & io_ex_datapathio_ex_Branch; // @[Datapath.scala 75:98:@846.4]
  assign _T_73 = 2'h2 == io_ex_datapathio_Forward_A; // @[Mux.scala 46:19:@850.4]
  assign _T_74 = _T_73 ? io_ex_datapathio_mem_alu_sum : io_ex_datapathio_ex_rs1_out; // @[Mux.scala 46:16:@851.4]
  assign _T_75 = 2'h1 == io_ex_datapathio_Forward_A; // @[Mux.scala 46:19:@852.4]
  assign _T_76 = _T_75 ? io_wb_datapathio_wb_reg_writedata : _T_74; // @[Mux.scala 46:16:@853.4]
  assign _T_77 = 2'h0 == io_ex_datapathio_Forward_A; // @[Mux.scala 46:19:@854.4]
  assign _T_79 = 2'h2 == io_ex_datapathio_Forward_B; // @[Mux.scala 46:19:@857.4]
  assign _T_80 = _T_79 ? io_ex_datapathio_mem_alu_sum : io_ex_datapathio_ex_rs2_out; // @[Mux.scala 46:16:@858.4]
  assign _T_81 = 2'h1 == io_ex_datapathio_Forward_B; // @[Mux.scala 46:19:@859.4]
  assign _T_82 = _T_81 ? io_wb_datapathio_wb_reg_writedata : _T_80; // @[Mux.scala 46:16:@860.4]
  assign _T_83 = 2'h0 == io_ex_datapathio_Forward_B; // @[Mux.scala 46:19:@861.4]
  assign operand_b = _T_83 ? io_ex_datapathio_ex_rs2_out : _T_82; // @[Mux.scala 46:16:@862.4]
  assign _T_86 = 3'h4 == io_wb_datapathio_wb_Mem_to_Reg; // @[Mux.scala 46:19:@867.4]
  assign _T_87 = _T_86 ? io_wb_datapathio_wb_aui_pc : io_wb_datapathio_wb_alu_sum; // @[Mux.scala 46:16:@868.4]
  assign _T_88 = 3'h3 == io_wb_datapathio_wb_Mem_to_Reg; // @[Mux.scala 46:19:@869.4]
  assign _T_89 = _T_88 ? io_wb_datapathio_wb_imm : _T_87; // @[Mux.scala 46:16:@870.4]
  assign _T_90 = 3'h2 == io_wb_datapathio_wb_Mem_to_Reg; // @[Mux.scala 46:19:@871.4]
  assign _T_91 = _T_90 ? io_wb_datapathio_wb_pc_4 : _T_89; // @[Mux.scala 46:16:@872.4]
  assign _T_92 = 3'h1 == io_wb_datapathio_wb_Mem_to_Reg; // @[Mux.scala 46:19:@873.4]
  assign _T_93 = _T_92 ? io_wb_datapathio_wb_dataout : _T_91; // @[Mux.scala 46:16:@874.4]
  assign _T_94 = 3'h0 == io_wb_datapathio_wb_Mem_to_Reg; // @[Mux.scala 46:19:@875.4]
  assign io_if_datapathio_if_new_pc = PC_Src ? ex_branch_addr : PC_4; // @[Datapath.scala 77:30:@849.4]
  assign io_if_datapathio_if_pc_4 = io_if_datapathio_if_pc + 32'h4; // @[Datapath.scala 67:28:@838.4]
  assign io_ex_datapathio_alu_b_src = io_ex_datapathio_ex_ALU_Src ? io_ex_datapathio_ex_imm : operand_b; // @[Datapath.scala 96:30:@865.4]
  assign io_ex_datapathio_ex_aui_pc = _T_60 + io_ex_datapathio_ex_imm; // @[Datapath.scala 72:30:@843.4]
  assign io_ex_datapathio_forward_rs2_out = _T_83 ? io_ex_datapathio_ex_rs2_out : _T_82; // @[Datapath.scala 98:36:@866.4]
  assign io_ex_datapathio_alu_a_src = _T_77 ? io_ex_datapathio_ex_rs1_out : _T_76; // @[Datapath.scala 81:30:@856.4]
  assign io_wb_datapathio_wb_reg_writedata = _T_94 ? io_wb_datapathio_wb_alu_sum : _T_93; // @[Datapath.scala 105:37:@877.4]
endmodule
module EX_MEM_Register( // @[:@879.2]
  input         clock, // @[:@880.4]
  input         reset, // @[:@881.4]
  input  [31:0] io_ex_alu_sum, // @[:@882.4]
  input  [31:0] io_ex_rs2_out, // @[:@882.4]
  input  [4:0]  io_ex_rd, // @[:@882.4]
  input  [31:0] io_ex_pc_4, // @[:@882.4]
  input  [31:0] io_ex_imm, // @[:@882.4]
  input  [31:0] io_ex_aui_pc, // @[:@882.4]
  input         io_ex_Mem_Read, // @[:@882.4]
  input         io_ex_Mem_Write, // @[:@882.4]
  input  [1:0]  io_ex_Data_Size, // @[:@882.4]
  input         io_ex_Load_Type, // @[:@882.4]
  input         io_ex_Reg_Write, // @[:@882.4]
  input  [2:0]  io_ex_Mem_to_Reg, // @[:@882.4]
  output        io_mem_Mem_Read, // @[:@882.4]
  output        io_mem_Mem_Write, // @[:@882.4]
  output [1:0]  io_mem_Data_Size, // @[:@882.4]
  output        io_mem_Load_Type, // @[:@882.4]
  output        io_mem_Reg_Write, // @[:@882.4]
  output [2:0]  io_mem_Mem_to_Reg, // @[:@882.4]
  output [31:0] io_mem_alu_sum, // @[:@882.4]
  output [31:0] io_mem_rs2_out, // @[:@882.4]
  output [4:0]  io_mem_rd, // @[:@882.4]
  output [31:0] io_mem_pc_4, // @[:@882.4]
  output [31:0] io_mem_imm, // @[:@882.4]
  output [31:0] io_mem_aui_pc // @[:@882.4]
);
  reg [31:0] alu_sum; // @[EX_MEM_Register.scala 53:30:@884.4]
  reg [31:0] _RAND_0;
  reg [31:0] rs2_out; // @[EX_MEM_Register.scala 54:30:@885.4]
  reg [31:0] _RAND_1;
  reg [4:0] rd; // @[EX_MEM_Register.scala 55:30:@886.4]
  reg [31:0] _RAND_2;
  reg [31:0] pc_4; // @[EX_MEM_Register.scala 56:30:@887.4]
  reg [31:0] _RAND_3;
  reg [31:0] imm; // @[EX_MEM_Register.scala 57:30:@888.4]
  reg [31:0] _RAND_4;
  reg [31:0] aui_pc; // @[EX_MEM_Register.scala 58:30:@889.4]
  reg [31:0] _RAND_5;
  reg  mem_read; // @[EX_MEM_Register.scala 60:30:@890.4]
  reg [31:0] _RAND_6;
  reg  mem_write; // @[EX_MEM_Register.scala 61:30:@891.4]
  reg [31:0] _RAND_7;
  reg [1:0] data_size; // @[EX_MEM_Register.scala 62:30:@892.4]
  reg [31:0] _RAND_8;
  reg  load_type; // @[EX_MEM_Register.scala 63:30:@893.4]
  reg [31:0] _RAND_9;
  reg  reg_write; // @[EX_MEM_Register.scala 64:30:@894.4]
  reg [31:0] _RAND_10;
  reg [2:0] mem_to_reg; // @[EX_MEM_Register.scala 65:30:@895.4]
  reg [31:0] _RAND_11;
  assign io_mem_Mem_Read = mem_read; // @[EX_MEM_Register.scala 88:23:@914.4]
  assign io_mem_Mem_Write = mem_write; // @[EX_MEM_Register.scala 89:23:@915.4]
  assign io_mem_Data_Size = data_size; // @[EX_MEM_Register.scala 90:23:@916.4]
  assign io_mem_Load_Type = load_type; // @[EX_MEM_Register.scala 91:23:@917.4]
  assign io_mem_Reg_Write = reg_write; // @[EX_MEM_Register.scala 92:23:@918.4]
  assign io_mem_Mem_to_Reg = mem_to_reg; // @[EX_MEM_Register.scala 93:23:@919.4]
  assign io_mem_alu_sum = alu_sum; // @[EX_MEM_Register.scala 82:23:@908.4]
  assign io_mem_rs2_out = rs2_out; // @[EX_MEM_Register.scala 83:23:@909.4]
  assign io_mem_rd = rd; // @[EX_MEM_Register.scala 84:23:@910.4]
  assign io_mem_pc_4 = pc_4; // @[EX_MEM_Register.scala 85:23:@911.4]
  assign io_mem_imm = imm; // @[EX_MEM_Register.scala 86:23:@912.4]
  assign io_mem_aui_pc = aui_pc; // @[EX_MEM_Register.scala 87:23:@913.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  alu_sum = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rs2_out = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rd = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  pc_4 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imm = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  aui_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_read = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_write = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  data_size = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  load_type = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_write = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_to_reg = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      alu_sum <= 32'h0;
    end else begin
      alu_sum <= io_ex_alu_sum;
    end
    if (reset) begin
      rs2_out <= 32'h0;
    end else begin
      rs2_out <= io_ex_rs2_out;
    end
    if (reset) begin
      rd <= 5'h0;
    end else begin
      rd <= io_ex_rd;
    end
    if (reset) begin
      pc_4 <= 32'h0;
    end else begin
      pc_4 <= io_ex_pc_4;
    end
    if (reset) begin
      imm <= 32'h0;
    end else begin
      imm <= io_ex_imm;
    end
    if (reset) begin
      aui_pc <= 32'h0;
    end else begin
      aui_pc <= io_ex_aui_pc;
    end
    if (reset) begin
      mem_read <= 1'h0;
    end else begin
      mem_read <= io_ex_Mem_Read;
    end
    if (reset) begin
      mem_write <= 1'h0;
    end else begin
      mem_write <= io_ex_Mem_Write;
    end
    if (reset) begin
      data_size <= 2'h0;
    end else begin
      data_size <= io_ex_Data_Size;
    end
    if (reset) begin
      load_type <= 1'h0;
    end else begin
      load_type <= io_ex_Load_Type;
    end
    if (reset) begin
      reg_write <= 1'h0;
    end else begin
      reg_write <= io_ex_Reg_Write;
    end
    if (reset) begin
      mem_to_reg <= 3'h0;
    end else begin
      mem_to_reg <= io_ex_Mem_to_Reg;
    end
  end
endmodule
module DataCache( // @[:@921.2]
  input         clock, // @[:@922.4]
  input  [31:0] io_addr, // @[:@924.4]
  input  [31:0] io_write_data, // @[:@924.4]
  input         io_Mem_Read, // @[:@924.4]
  input         io_Mem_Write, // @[:@924.4]
  input  [1:0]  io_Data_Size, // @[:@924.4]
  input         io_Load_Type, // @[:@924.4]
  output [31:0] io_data_out // @[:@924.4]
);
  reg [31:0] cache [0:31]; // @[DataCache.scala 41:18:@926.4]
  reg [31:0] _RAND_0;
  wire [31:0] cache__T_35_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_35_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_37_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_37_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_39_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_39_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_42_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_42_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_51_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_51_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_54_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_54_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_75_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_75_addr; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] cache__T_72_data; // @[DataCache.scala 41:18:@926.4]
  wire [4:0] cache__T_72_addr; // @[DataCache.scala 41:18:@926.4]
  wire  cache__T_72_mask; // @[DataCache.scala 41:18:@926.4]
  wire  cache__T_72_en; // @[DataCache.scala 41:18:@926.4]
  wire [31:0] fix_addr; // @[DataCache.scala 44:26:@927.4]
  wire [15:0] _T_23; // @[DataCache.scala 48:48:@928.4]
  wire [31:0] _T_24; // @[Cat.scala 30:58:@929.4]
  wire [7:0] _T_26; // @[DataCache.scala 49:48:@930.4]
  wire [31:0] _T_27; // @[Cat.scala 30:58:@931.4]
  wire  _T_28; // @[Mux.scala 46:19:@932.4]
  wire [31:0] _T_29; // @[Mux.scala 46:16:@933.4]
  wire  _T_30; // @[Mux.scala 46:19:@934.4]
  wire [31:0] _T_31; // @[Mux.scala 46:16:@935.4]
  wire  _T_32; // @[Mux.scala 46:19:@936.4]
  wire [31:0] write_data; // @[Mux.scala 46:16:@937.4]
  wire [2:0] _T_33; // @[Cat.scala 30:58:@938.4]
  wire [15:0] _T_40; // @[DataCache.scala 54:38:@945.4]
  wire [15:0] _T_43; // @[DataCache.scala 55:40:@948.4]
  wire [15:0] _T_44; // @[DataCache.scala 55:54:@949.4]
  wire [46:0] _GEN_18; // @[DataCache.scala 55:57:@950.4]
  wire [46:0] _T_46; // @[DataCache.scala 55:57:@950.4]
  wire [46:0] _T_48; // @[DataCache.scala 55:66:@951.4]
  wire [46:0] _T_49; // @[DataCache.scala 55:81:@952.4]
  wire [7:0] _T_52; // @[DataCache.scala 56:38:@955.4]
  wire [7:0] _T_55; // @[DataCache.scala 57:40:@958.4]
  wire [7:0] _T_56; // @[DataCache.scala 57:53:@959.4]
  wire [38:0] _GEN_19; // @[DataCache.scala 57:56:@960.4]
  wire [38:0] _T_58; // @[DataCache.scala 57:56:@960.4]
  wire [38:0] _T_60; // @[DataCache.scala 57:65:@961.4]
  wire [38:0] _T_61; // @[DataCache.scala 57:80:@962.4]
  wire  _T_62; // @[Mux.scala 46:19:@963.4]
  wire [38:0] _T_63; // @[Mux.scala 46:16:@964.4]
  wire  _T_64; // @[Mux.scala 46:19:@965.4]
  wire [38:0] _T_65; // @[Mux.scala 46:16:@966.4]
  wire  _T_66; // @[Mux.scala 46:19:@967.4]
  wire [46:0] _T_67; // @[Mux.scala 46:16:@968.4]
  wire  _T_68; // @[Mux.scala 46:19:@969.4]
  wire [46:0] _T_69; // @[Mux.scala 46:16:@970.4]
  wire  _T_70; // @[Mux.scala 46:19:@971.4]
  wire [46:0] read_data; // @[Mux.scala 46:16:@972.4]
  wire [46:0] _T_79; // @[DataCache.scala 61:21:@981.4]
  assign cache__T_35_addr = fix_addr[4:0];
  assign cache__T_35_data = cache[cache__T_35_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_37_addr = fix_addr[4:0];
  assign cache__T_37_data = cache[cache__T_37_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_39_addr = fix_addr[4:0];
  assign cache__T_39_data = cache[cache__T_39_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_42_addr = fix_addr[4:0];
  assign cache__T_42_data = cache[cache__T_42_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_51_addr = fix_addr[4:0];
  assign cache__T_51_data = cache[cache__T_51_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_54_addr = fix_addr[4:0];
  assign cache__T_54_data = cache[cache__T_54_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_75_addr = fix_addr[4:0];
  assign cache__T_75_data = cache[cache__T_75_addr]; // @[DataCache.scala 41:18:@926.4]
  assign cache__T_72_data = io_Mem_Write ? write_data : cache__T_75_data;
  assign cache__T_72_addr = fix_addr[4:0];
  assign cache__T_72_mask = 1'h1;
  assign cache__T_72_en = 1'h1;
  assign fix_addr = io_addr / 32'h4; // @[DataCache.scala 44:26:@927.4]
  assign _T_23 = io_write_data[15:0]; // @[DataCache.scala 48:48:@928.4]
  assign _T_24 = {16'h0,_T_23}; // @[Cat.scala 30:58:@929.4]
  assign _T_26 = io_write_data[7:0]; // @[DataCache.scala 49:48:@930.4]
  assign _T_27 = {24'h0,_T_26}; // @[Cat.scala 30:58:@931.4]
  assign _T_28 = 2'h2 == io_Data_Size; // @[Mux.scala 46:19:@932.4]
  assign _T_29 = _T_28 ? _T_27 : io_write_data; // @[Mux.scala 46:16:@933.4]
  assign _T_30 = 2'h1 == io_Data_Size; // @[Mux.scala 46:19:@934.4]
  assign _T_31 = _T_30 ? _T_24 : _T_29; // @[Mux.scala 46:16:@935.4]
  assign _T_32 = 2'h0 == io_Data_Size; // @[Mux.scala 46:19:@936.4]
  assign write_data = _T_32 ? io_write_data : _T_31; // @[Mux.scala 46:16:@937.4]
  assign _T_33 = {io_Data_Size,io_Load_Type}; // @[Cat.scala 30:58:@938.4]
  assign _T_40 = cache__T_39_data[15:0]; // @[DataCache.scala 54:38:@945.4]
  assign _T_43 = cache__T_42_data[15:0]; // @[DataCache.scala 55:40:@948.4]
  assign _T_44 = $signed(_T_43); // @[DataCache.scala 55:54:@949.4]
  assign _GEN_18 = {{31{_T_44[15]}},_T_44}; // @[DataCache.scala 55:57:@950.4]
  assign _T_46 = $signed(_GEN_18) << 5'h10; // @[DataCache.scala 55:57:@950.4]
  assign _T_48 = $signed(_T_46) >>> 5'h10; // @[DataCache.scala 55:66:@951.4]
  assign _T_49 = $unsigned(_T_48); // @[DataCache.scala 55:81:@952.4]
  assign _T_52 = cache__T_51_data[7:0]; // @[DataCache.scala 56:38:@955.4]
  assign _T_55 = cache__T_54_data[7:0]; // @[DataCache.scala 57:40:@958.4]
  assign _T_56 = $signed(_T_55); // @[DataCache.scala 57:53:@959.4]
  assign _GEN_19 = {{31{_T_56[7]}},_T_56}; // @[DataCache.scala 57:56:@960.4]
  assign _T_58 = $signed(_GEN_19) << 5'h18; // @[DataCache.scala 57:56:@960.4]
  assign _T_60 = $signed(_T_58) >>> 5'h18; // @[DataCache.scala 57:65:@961.4]
  assign _T_61 = $unsigned(_T_60); // @[DataCache.scala 57:80:@962.4]
  assign _T_62 = 3'h4 == _T_33; // @[Mux.scala 46:19:@963.4]
  assign _T_63 = _T_62 ? _T_61 : {{7'd0}, cache__T_35_data}; // @[Mux.scala 46:16:@964.4]
  assign _T_64 = 3'h5 == _T_33; // @[Mux.scala 46:19:@965.4]
  assign _T_65 = _T_64 ? {{31'd0}, _T_52} : _T_63; // @[Mux.scala 46:16:@966.4]
  assign _T_66 = 3'h2 == _T_33; // @[Mux.scala 46:19:@967.4]
  assign _T_67 = _T_66 ? _T_49 : {{8'd0}, _T_65}; // @[Mux.scala 46:16:@968.4]
  assign _T_68 = 3'h3 == _T_33; // @[Mux.scala 46:19:@969.4]
  assign _T_69 = _T_68 ? {{31'd0}, _T_40} : _T_67; // @[Mux.scala 46:16:@970.4]
  assign _T_70 = 3'h1 == _T_33; // @[Mux.scala 46:19:@971.4]
  assign read_data = _T_70 ? {{15'd0}, cache__T_37_data} : _T_69; // @[Mux.scala 46:16:@972.4]
  assign _T_79 = io_Mem_Read ? read_data : 47'h0; // @[DataCache.scala 61:21:@981.4]
  assign io_data_out = _T_79[31:0]; // @[DataCache.scala 61:15:@982.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    cache[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(cache__T_72_en & cache__T_72_mask) begin
      cache[cache__T_72_addr] <= cache__T_72_data; // @[DataCache.scala 41:18:@926.4]
    end
  end
endmodule
module MEM_WB_Register( // @[:@984.2]
  input         clock, // @[:@985.4]
  input         reset, // @[:@986.4]
  input  [31:0] io_mem_dataout, // @[:@987.4]
  input  [31:0] io_mem_alu_sum, // @[:@987.4]
  input  [4:0]  io_mem_rd, // @[:@987.4]
  input  [31:0] io_mem_pc_4, // @[:@987.4]
  input  [31:0] io_mem_imm, // @[:@987.4]
  input  [31:0] io_mem_aui_pc, // @[:@987.4]
  input  [2:0]  io_mem_Mem_to_Reg, // @[:@987.4]
  input         io_mem_Reg_Write, // @[:@987.4]
  output [2:0]  io_wb_Mem_to_Reg, // @[:@987.4]
  output        io_wb_Reg_Write, // @[:@987.4]
  output [31:0] io_wb_dataout, // @[:@987.4]
  output [31:0] io_wb_alu_sum, // @[:@987.4]
  output [4:0]  io_wb_rd, // @[:@987.4]
  output [31:0] io_wb_pc_4, // @[:@987.4]
  output [31:0] io_wb_imm, // @[:@987.4]
  output [31:0] io_wb_aui_pc // @[:@987.4]
);
  reg [31:0] dataout; // @[MEM_WB_Register.scala 43:28:@989.4]
  reg [31:0] _RAND_0;
  reg [31:0] alu_sum; // @[MEM_WB_Register.scala 44:28:@990.4]
  reg [31:0] _RAND_1;
  reg [4:0] rd; // @[MEM_WB_Register.scala 45:28:@991.4]
  reg [31:0] _RAND_2;
  reg [31:0] pc_4; // @[MEM_WB_Register.scala 46:28:@992.4]
  reg [31:0] _RAND_3;
  reg [31:0] imm; // @[MEM_WB_Register.scala 47:28:@993.4]
  reg [31:0] _RAND_4;
  reg [31:0] aui_pc; // @[MEM_WB_Register.scala 48:28:@994.4]
  reg [31:0] _RAND_5;
  reg [2:0] mem_to_reg; // @[MEM_WB_Register.scala 49:28:@995.4]
  reg [31:0] _RAND_6;
  reg  reg_write; // @[MEM_WB_Register.scala 50:28:@996.4]
  reg [31:0] _RAND_7;
  assign io_wb_Mem_to_Reg = mem_to_reg; // @[MEM_WB_Register.scala 63:21:@1005.4]
  assign io_wb_Reg_Write = reg_write; // @[MEM_WB_Register.scala 64:21:@1006.4]
  assign io_wb_dataout = dataout; // @[MEM_WB_Register.scala 65:21:@1007.4]
  assign io_wb_alu_sum = alu_sum; // @[MEM_WB_Register.scala 66:21:@1008.4]
  assign io_wb_rd = rd; // @[MEM_WB_Register.scala 67:21:@1009.4]
  assign io_wb_pc_4 = pc_4; // @[MEM_WB_Register.scala 68:21:@1010.4]
  assign io_wb_imm = imm; // @[MEM_WB_Register.scala 69:21:@1011.4]
  assign io_wb_aui_pc = aui_pc; // @[MEM_WB_Register.scala 70:21:@1012.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dataout = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  alu_sum = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rd = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  pc_4 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imm = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  aui_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_to_reg = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_write = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      dataout <= 32'h0;
    end else begin
      dataout <= io_mem_dataout;
    end
    if (reset) begin
      alu_sum <= 32'h0;
    end else begin
      alu_sum <= io_mem_alu_sum;
    end
    if (reset) begin
      rd <= 5'h0;
    end else begin
      rd <= io_mem_rd;
    end
    if (reset) begin
      pc_4 <= 32'h0;
    end else begin
      pc_4 <= io_mem_pc_4;
    end
    if (reset) begin
      imm <= 32'h0;
    end else begin
      imm <= io_mem_imm;
    end
    if (reset) begin
      aui_pc <= 32'h0;
    end else begin
      aui_pc <= io_mem_aui_pc;
    end
    if (reset) begin
      mem_to_reg <= 3'h0;
    end else begin
      mem_to_reg <= io_mem_Mem_to_Reg;
    end
    if (reset) begin
      reg_write <= 1'h0;
    end else begin
      reg_write <= io_mem_Reg_Write;
    end
  end
endmodule
module Forward( // @[:@1014.2]
  input        io_ex_mem_Reg_Write, // @[:@1017.4]
  input  [4:0] io_ex_mem_rd, // @[:@1017.4]
  input        io_mem_wb_Reg_Write, // @[:@1017.4]
  input  [4:0] io_mem_wb_rd, // @[:@1017.4]
  input  [4:0] io_id_ex_rs1, // @[:@1017.4]
  input  [4:0] io_id_ex_rs2, // @[:@1017.4]
  output [1:0] io_Forward_A, // @[:@1017.4]
  output [1:0] io_Forward_B // @[:@1017.4]
);
  wire  _T_23; // @[Forward.scala 43:35:@1020.4]
  wire  _T_24; // @[Forward.scala 42:51:@1021.4]
  wire  _T_25; // @[Forward.scala 44:36:@1022.4]
  wire  ex_mem_a_con; // @[Forward.scala 43:51:@1023.4]
  wire  _T_28; // @[Forward.scala 46:35:@1025.4]
  wire  _T_29; // @[Forward.scala 45:51:@1026.4]
  wire  _T_31; // @[Forward.scala 47:22:@1027.4]
  wire  _T_32; // @[Forward.scala 46:51:@1028.4]
  wire  _T_33; // @[Forward.scala 48:36:@1029.4]
  wire  ex_wb_a_con; // @[Forward.scala 47:51:@1030.4]
  wire  _T_38; // @[Forward.scala 51:36:@1034.4]
  wire  ex_mem_b_con; // @[Forward.scala 50:51:@1035.4]
  wire  _T_44; // @[Forward.scala 54:22:@1039.4]
  wire  _T_45; // @[Forward.scala 53:51:@1040.4]
  wire  _T_46; // @[Forward.scala 55:36:@1041.4]
  wire  ex_wb_b_con; // @[Forward.scala 54:51:@1042.4]
  assign _T_23 = io_ex_mem_rd != 5'h0; // @[Forward.scala 43:35:@1020.4]
  assign _T_24 = io_ex_mem_Reg_Write & _T_23; // @[Forward.scala 42:51:@1021.4]
  assign _T_25 = io_ex_mem_rd == io_id_ex_rs1; // @[Forward.scala 44:36:@1022.4]
  assign ex_mem_a_con = _T_24 & _T_25; // @[Forward.scala 43:51:@1023.4]
  assign _T_28 = io_mem_wb_rd != 5'h0; // @[Forward.scala 46:35:@1025.4]
  assign _T_29 = io_mem_wb_Reg_Write & _T_28; // @[Forward.scala 45:51:@1026.4]
  assign _T_31 = ex_mem_a_con == 1'h0; // @[Forward.scala 47:22:@1027.4]
  assign _T_32 = _T_29 & _T_31; // @[Forward.scala 46:51:@1028.4]
  assign _T_33 = io_mem_wb_rd == io_id_ex_rs1; // @[Forward.scala 48:36:@1029.4]
  assign ex_wb_a_con = _T_32 & _T_33; // @[Forward.scala 47:51:@1030.4]
  assign _T_38 = io_ex_mem_rd == io_id_ex_rs2; // @[Forward.scala 51:36:@1034.4]
  assign ex_mem_b_con = _T_24 & _T_38; // @[Forward.scala 50:51:@1035.4]
  assign _T_44 = ex_mem_b_con == 1'h0; // @[Forward.scala 54:22:@1039.4]
  assign _T_45 = _T_29 & _T_44; // @[Forward.scala 53:51:@1040.4]
  assign _T_46 = io_mem_wb_rd == io_id_ex_rs2; // @[Forward.scala 55:36:@1041.4]
  assign ex_wb_b_con = _T_45 & _T_46; // @[Forward.scala 54:51:@1042.4]
  assign io_Forward_A = {ex_mem_a_con,ex_wb_a_con}; // @[Forward.scala 57:16:@1044.4]
  assign io_Forward_B = {ex_mem_b_con,ex_wb_b_con}; // @[Forward.scala 58:16:@1046.4]
endmodule
module Tile( // @[:@1048.2]
  input         clock, // @[:@1049.4]
  input         reset, // @[:@1050.4]
  input         io_pc_write, // @[:@1051.4]
  input         io_if_id_write, // @[:@1051.4]
  input         io_if_flush, // @[:@1051.4]
  output [31:0] io_if_pc_out, // @[:@1051.4]
  output [31:0] io_if_next_pc, // @[:@1051.4]
  output [4:0]  io_id_rs1, // @[:@1051.4]
  output [4:0]  io_id_rs2, // @[:@1051.4]
  output [31:0] io_id_rs1_out, // @[:@1051.4]
  output [31:0] io_id_rs2_out, // @[:@1051.4]
  output [31:0] io_ex_rs1_out, // @[:@1051.4]
  output [31:0] io_ex_rs2_out, // @[:@1051.4]
  output [31:0] io_ex_alu_sum, // @[:@1051.4]
  output        io_ex_alu_conflag, // @[:@1051.4]
  output [4:0]  io_ex_rd, // @[:@1051.4]
  output [4:0]  io_mem_rd, // @[:@1051.4]
  output [31:0] io_mem_alu_sum, // @[:@1051.4]
  output [31:0] io_mem_writedata, // @[:@1051.4]
  output [31:0] io_mem_dataout, // @[:@1051.4]
  output [4:0]  io_wb_rd, // @[:@1051.4]
  output [31:0] io_wb_registerwrite, // @[:@1051.4]
  output [1:0]  io_Forward_A, // @[:@1051.4]
  output [1:0]  io_Forward_B // @[:@1051.4]
);
  wire  pc_clock; // @[Tile.scala 50:31:@1053.4]
  wire  pc_reset; // @[Tile.scala 50:31:@1053.4]
  wire [31:0] pc_io_addr_input; // @[Tile.scala 50:31:@1053.4]
  wire  pc_io_pc_write; // @[Tile.scala 50:31:@1053.4]
  wire [31:0] pc_io_pc_out; // @[Tile.scala 50:31:@1053.4]
  wire  instcache_clock; // @[Tile.scala 51:31:@1056.4]
  wire [31:0] instcache_io_addr; // @[Tile.scala 51:31:@1056.4]
  wire [31:0] instcache_io_inst; // @[Tile.scala 51:31:@1056.4]
  wire  if_id_register_clock; // @[Tile.scala 52:31:@1059.4]
  wire  if_id_register_reset; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_if_pc; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_if_inst; // @[Tile.scala 52:31:@1059.4]
  wire  if_id_register_io_if_id_write; // @[Tile.scala 52:31:@1059.4]
  wire  if_id_register_io_if_flush; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_if_pc_4; // @[Tile.scala 52:31:@1059.4]
  wire [4:0] if_id_register_io_id_rs1; // @[Tile.scala 52:31:@1059.4]
  wire [4:0] if_id_register_io_id_rs2; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_id_pc; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_id_pc_4; // @[Tile.scala 52:31:@1059.4]
  wire [31:0] if_id_register_io_id_inst; // @[Tile.scala 52:31:@1059.4]
  wire  regfile_clock; // @[Tile.scala 53:31:@1062.4]
  wire [4:0] regfile_io_rs1; // @[Tile.scala 53:31:@1062.4]
  wire [4:0] regfile_io_rs2; // @[Tile.scala 53:31:@1062.4]
  wire [4:0] regfile_io_rd; // @[Tile.scala 53:31:@1062.4]
  wire [31:0] regfile_io_wdata; // @[Tile.scala 53:31:@1062.4]
  wire  regfile_io_regwrite; // @[Tile.scala 53:31:@1062.4]
  wire [31:0] regfile_io_rs1_out; // @[Tile.scala 53:31:@1062.4]
  wire [31:0] regfile_io_rs2_out; // @[Tile.scala 53:31:@1062.4]
  wire [31:0] immgen_io_inst_in; // @[Tile.scala 54:31:@1065.4]
  wire [2:0] immgen_io_imm_sel; // @[Tile.scala 54:31:@1065.4]
  wire [31:0] immgen_io_imm; // @[Tile.scala 54:31:@1065.4]
  wire [31:0] control_io_inst; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Reg_Write; // @[Tile.scala 55:31:@1068.4]
  wire [2:0] control_io_Imm_Sel; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_ALU_Src; // @[Tile.scala 55:31:@1068.4]
  wire [4:0] control_io_ALUOp; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Branch; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Branch_Src; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Mem_Read; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Mem_Write; // @[Tile.scala 55:31:@1068.4]
  wire [1:0] control_io_Data_Size; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Load_Type; // @[Tile.scala 55:31:@1068.4]
  wire [2:0] control_io_Mem_to_Reg; // @[Tile.scala 55:31:@1068.4]
  wire  control_io_Jump_Type; // @[Tile.scala 55:31:@1068.4]
  wire  id_ex_register_clock; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_reset; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_pc; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_pc_4; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_rs1_out; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_rs2_out; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_imm; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_id_inst; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_id_rs1; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_id_rs2; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ALU_Src; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_ALUOp; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Branch; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Branch_Src; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Jump_Type; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Mem_Read; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Mem_Write; // @[Tile.scala 56:31:@1071.4]
  wire [1:0] id_ex_register_io_Data_Size; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Load_Type; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_Reg_Write; // @[Tile.scala 56:31:@1071.4]
  wire [2:0] id_ex_register_io_Mem_to_Reg; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_ALU_Src; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_ex_ALUOp; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Branch; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Branch_Src; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Jump_Type; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Mem_Read; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Mem_Write; // @[Tile.scala 56:31:@1071.4]
  wire [1:0] id_ex_register_io_ex_Data_Size; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Load_Type; // @[Tile.scala 56:31:@1071.4]
  wire  id_ex_register_io_ex_Reg_Write; // @[Tile.scala 56:31:@1071.4]
  wire [2:0] id_ex_register_io_ex_Mem_to_Reg; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_ex_pc; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_ex_pc_4; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_ex_rs1_out; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_ex_rs2_out; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_ex_rd; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] id_ex_register_io_ex_imm; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_ex_rs1; // @[Tile.scala 56:31:@1071.4]
  wire [4:0] id_ex_register_io_ex_rs2; // @[Tile.scala 56:31:@1071.4]
  wire [31:0] alu_io_Src_A; // @[Tile.scala 57:31:@1074.4]
  wire [31:0] alu_io_Src_B; // @[Tile.scala 57:31:@1074.4]
  wire [4:0] alu_io_ALUOp; // @[Tile.scala 57:31:@1074.4]
  wire [31:0] alu_io_Sum; // @[Tile.scala 57:31:@1074.4]
  wire  alu_io_Conflag; // @[Tile.scala 57:31:@1074.4]
  wire [31:0] datapath_io_if_datapathio_if_pc; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_if_datapathio_if_new_pc; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_if_datapathio_if_pc_4; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_ex_rs1_out; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_ex_rs2_out; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_ex_imm; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_ex_pc; // @[Tile.scala 58:31:@1077.4]
  wire  datapath_io_ex_datapathio_ex_ALU_Src; // @[Tile.scala 58:31:@1077.4]
  wire  datapath_io_ex_datapathio_ex_Branch; // @[Tile.scala 58:31:@1077.4]
  wire  datapath_io_ex_datapathio_ex_alu_conflag; // @[Tile.scala 58:31:@1077.4]
  wire  datapath_io_ex_datapathio_ex_Branch_Src; // @[Tile.scala 58:31:@1077.4]
  wire  datapath_io_ex_datapathio_ex_Jump_Type; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_mem_alu_sum; // @[Tile.scala 58:31:@1077.4]
  wire [1:0] datapath_io_ex_datapathio_Forward_A; // @[Tile.scala 58:31:@1077.4]
  wire [1:0] datapath_io_ex_datapathio_Forward_B; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_alu_b_src; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_ex_aui_pc; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_forward_rs2_out; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_ex_datapathio_alu_a_src; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_alu_sum; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_dataout; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_pc_4; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_imm; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_aui_pc; // @[Tile.scala 58:31:@1077.4]
  wire [2:0] datapath_io_wb_datapathio_wb_Mem_to_Reg; // @[Tile.scala 58:31:@1077.4]
  wire [31:0] datapath_io_wb_datapathio_wb_reg_writedata; // @[Tile.scala 58:31:@1077.4]
  wire  ex_mem_register_clock; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_reset; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_ex_alu_sum; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_ex_rs2_out; // @[Tile.scala 59:31:@1080.4]
  wire [4:0] ex_mem_register_io_ex_rd; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_ex_pc_4; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_ex_imm; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_ex_aui_pc; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_ex_Mem_Read; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_ex_Mem_Write; // @[Tile.scala 59:31:@1080.4]
  wire [1:0] ex_mem_register_io_ex_Data_Size; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_ex_Load_Type; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_ex_Reg_Write; // @[Tile.scala 59:31:@1080.4]
  wire [2:0] ex_mem_register_io_ex_Mem_to_Reg; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_mem_Mem_Read; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_mem_Mem_Write; // @[Tile.scala 59:31:@1080.4]
  wire [1:0] ex_mem_register_io_mem_Data_Size; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_mem_Load_Type; // @[Tile.scala 59:31:@1080.4]
  wire  ex_mem_register_io_mem_Reg_Write; // @[Tile.scala 59:31:@1080.4]
  wire [2:0] ex_mem_register_io_mem_Mem_to_Reg; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_mem_alu_sum; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_mem_rs2_out; // @[Tile.scala 59:31:@1080.4]
  wire [4:0] ex_mem_register_io_mem_rd; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_mem_pc_4; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_mem_imm; // @[Tile.scala 59:31:@1080.4]
  wire [31:0] ex_mem_register_io_mem_aui_pc; // @[Tile.scala 59:31:@1080.4]
  wire  datacache_clock; // @[Tile.scala 60:31:@1083.4]
  wire [31:0] datacache_io_addr; // @[Tile.scala 60:31:@1083.4]
  wire [31:0] datacache_io_write_data; // @[Tile.scala 60:31:@1083.4]
  wire  datacache_io_Mem_Read; // @[Tile.scala 60:31:@1083.4]
  wire  datacache_io_Mem_Write; // @[Tile.scala 60:31:@1083.4]
  wire [1:0] datacache_io_Data_Size; // @[Tile.scala 60:31:@1083.4]
  wire  datacache_io_Load_Type; // @[Tile.scala 60:31:@1083.4]
  wire [31:0] datacache_io_data_out; // @[Tile.scala 60:31:@1083.4]
  wire  mem_wb_register_clock; // @[Tile.scala 61:31:@1086.4]
  wire  mem_wb_register_reset; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_mem_dataout; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_mem_alu_sum; // @[Tile.scala 61:31:@1086.4]
  wire [4:0] mem_wb_register_io_mem_rd; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_mem_pc_4; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_mem_imm; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_mem_aui_pc; // @[Tile.scala 61:31:@1086.4]
  wire [2:0] mem_wb_register_io_mem_Mem_to_Reg; // @[Tile.scala 61:31:@1086.4]
  wire  mem_wb_register_io_mem_Reg_Write; // @[Tile.scala 61:31:@1086.4]
  wire [2:0] mem_wb_register_io_wb_Mem_to_Reg; // @[Tile.scala 61:31:@1086.4]
  wire  mem_wb_register_io_wb_Reg_Write; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_wb_dataout; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_wb_alu_sum; // @[Tile.scala 61:31:@1086.4]
  wire [4:0] mem_wb_register_io_wb_rd; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_wb_pc_4; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_wb_imm; // @[Tile.scala 61:31:@1086.4]
  wire [31:0] mem_wb_register_io_wb_aui_pc; // @[Tile.scala 61:31:@1086.4]
  wire  forward_io_ex_mem_Reg_Write; // @[Tile.scala 62:31:@1089.4]
  wire [4:0] forward_io_ex_mem_rd; // @[Tile.scala 62:31:@1089.4]
  wire  forward_io_mem_wb_Reg_Write; // @[Tile.scala 62:31:@1089.4]
  wire [4:0] forward_io_mem_wb_rd; // @[Tile.scala 62:31:@1089.4]
  wire [4:0] forward_io_id_ex_rs1; // @[Tile.scala 62:31:@1089.4]
  wire [4:0] forward_io_id_ex_rs2; // @[Tile.scala 62:31:@1089.4]
  wire [1:0] forward_io_Forward_A; // @[Tile.scala 62:31:@1089.4]
  wire [1:0] forward_io_Forward_B; // @[Tile.scala 62:31:@1089.4]
  PC pc ( // @[Tile.scala 50:31:@1053.4]
    .clock(pc_clock),
    .reset(pc_reset),
    .io_addr_input(pc_io_addr_input),
    .io_pc_write(pc_io_pc_write),
    .io_pc_out(pc_io_pc_out)
  );
  InstCache instcache ( // @[Tile.scala 51:31:@1056.4]
    .clock(instcache_clock),
    .io_addr(instcache_io_addr),
    .io_inst(instcache_io_inst)
  );
  IF_ID_Register if_id_register ( // @[Tile.scala 52:31:@1059.4]
    .clock(if_id_register_clock),
    .reset(if_id_register_reset),
    .io_if_pc(if_id_register_io_if_pc),
    .io_if_inst(if_id_register_io_if_inst),
    .io_if_id_write(if_id_register_io_if_id_write),
    .io_if_flush(if_id_register_io_if_flush),
    .io_if_pc_4(if_id_register_io_if_pc_4),
    .io_id_rs1(if_id_register_io_id_rs1),
    .io_id_rs2(if_id_register_io_id_rs2),
    .io_id_pc(if_id_register_io_id_pc),
    .io_id_pc_4(if_id_register_io_id_pc_4),
    .io_id_inst(if_id_register_io_id_inst)
  );
  RegFile regfile ( // @[Tile.scala 53:31:@1062.4]
    .clock(regfile_clock),
    .io_rs1(regfile_io_rs1),
    .io_rs2(regfile_io_rs2),
    .io_rd(regfile_io_rd),
    .io_wdata(regfile_io_wdata),
    .io_regwrite(regfile_io_regwrite),
    .io_rs1_out(regfile_io_rs1_out),
    .io_rs2_out(regfile_io_rs2_out)
  );
  ImmGen immgen ( // @[Tile.scala 54:31:@1065.4]
    .io_inst_in(immgen_io_inst_in),
    .io_imm_sel(immgen_io_imm_sel),
    .io_imm(immgen_io_imm)
  );
  Control control ( // @[Tile.scala 55:31:@1068.4]
    .io_inst(control_io_inst),
    .io_Reg_Write(control_io_Reg_Write),
    .io_Imm_Sel(control_io_Imm_Sel),
    .io_ALU_Src(control_io_ALU_Src),
    .io_ALUOp(control_io_ALUOp),
    .io_Branch(control_io_Branch),
    .io_Branch_Src(control_io_Branch_Src),
    .io_Mem_Read(control_io_Mem_Read),
    .io_Mem_Write(control_io_Mem_Write),
    .io_Data_Size(control_io_Data_Size),
    .io_Load_Type(control_io_Load_Type),
    .io_Mem_to_Reg(control_io_Mem_to_Reg),
    .io_Jump_Type(control_io_Jump_Type)
  );
  ID_EX_Register id_ex_register ( // @[Tile.scala 56:31:@1071.4]
    .clock(id_ex_register_clock),
    .reset(id_ex_register_reset),
    .io_id_pc(id_ex_register_io_id_pc),
    .io_id_pc_4(id_ex_register_io_id_pc_4),
    .io_id_rs1_out(id_ex_register_io_id_rs1_out),
    .io_id_rs2_out(id_ex_register_io_id_rs2_out),
    .io_id_imm(id_ex_register_io_id_imm),
    .io_id_inst(id_ex_register_io_id_inst),
    .io_id_rs1(id_ex_register_io_id_rs1),
    .io_id_rs2(id_ex_register_io_id_rs2),
    .io_ALU_Src(id_ex_register_io_ALU_Src),
    .io_ALUOp(id_ex_register_io_ALUOp),
    .io_Branch(id_ex_register_io_Branch),
    .io_Branch_Src(id_ex_register_io_Branch_Src),
    .io_Jump_Type(id_ex_register_io_Jump_Type),
    .io_Mem_Read(id_ex_register_io_Mem_Read),
    .io_Mem_Write(id_ex_register_io_Mem_Write),
    .io_Data_Size(id_ex_register_io_Data_Size),
    .io_Load_Type(id_ex_register_io_Load_Type),
    .io_Reg_Write(id_ex_register_io_Reg_Write),
    .io_Mem_to_Reg(id_ex_register_io_Mem_to_Reg),
    .io_ex_ALU_Src(id_ex_register_io_ex_ALU_Src),
    .io_ex_ALUOp(id_ex_register_io_ex_ALUOp),
    .io_ex_Branch(id_ex_register_io_ex_Branch),
    .io_ex_Branch_Src(id_ex_register_io_ex_Branch_Src),
    .io_ex_Jump_Type(id_ex_register_io_ex_Jump_Type),
    .io_ex_Mem_Read(id_ex_register_io_ex_Mem_Read),
    .io_ex_Mem_Write(id_ex_register_io_ex_Mem_Write),
    .io_ex_Data_Size(id_ex_register_io_ex_Data_Size),
    .io_ex_Load_Type(id_ex_register_io_ex_Load_Type),
    .io_ex_Reg_Write(id_ex_register_io_ex_Reg_Write),
    .io_ex_Mem_to_Reg(id_ex_register_io_ex_Mem_to_Reg),
    .io_ex_pc(id_ex_register_io_ex_pc),
    .io_ex_pc_4(id_ex_register_io_ex_pc_4),
    .io_ex_rs1_out(id_ex_register_io_ex_rs1_out),
    .io_ex_rs2_out(id_ex_register_io_ex_rs2_out),
    .io_ex_rd(id_ex_register_io_ex_rd),
    .io_ex_imm(id_ex_register_io_ex_imm),
    .io_ex_rs1(id_ex_register_io_ex_rs1),
    .io_ex_rs2(id_ex_register_io_ex_rs2)
  );
  ALU alu ( // @[Tile.scala 57:31:@1074.4]
    .io_Src_A(alu_io_Src_A),
    .io_Src_B(alu_io_Src_B),
    .io_ALUOp(alu_io_ALUOp),
    .io_Sum(alu_io_Sum),
    .io_Conflag(alu_io_Conflag)
  );
  Datapath datapath ( // @[Tile.scala 58:31:@1077.4]
    .io_if_datapathio_if_pc(datapath_io_if_datapathio_if_pc),
    .io_if_datapathio_if_new_pc(datapath_io_if_datapathio_if_new_pc),
    .io_if_datapathio_if_pc_4(datapath_io_if_datapathio_if_pc_4),
    .io_ex_datapathio_ex_rs1_out(datapath_io_ex_datapathio_ex_rs1_out),
    .io_ex_datapathio_ex_rs2_out(datapath_io_ex_datapathio_ex_rs2_out),
    .io_ex_datapathio_ex_imm(datapath_io_ex_datapathio_ex_imm),
    .io_ex_datapathio_ex_pc(datapath_io_ex_datapathio_ex_pc),
    .io_ex_datapathio_ex_ALU_Src(datapath_io_ex_datapathio_ex_ALU_Src),
    .io_ex_datapathio_ex_Branch(datapath_io_ex_datapathio_ex_Branch),
    .io_ex_datapathio_ex_alu_conflag(datapath_io_ex_datapathio_ex_alu_conflag),
    .io_ex_datapathio_ex_Branch_Src(datapath_io_ex_datapathio_ex_Branch_Src),
    .io_ex_datapathio_ex_Jump_Type(datapath_io_ex_datapathio_ex_Jump_Type),
    .io_ex_datapathio_mem_alu_sum(datapath_io_ex_datapathio_mem_alu_sum),
    .io_ex_datapathio_Forward_A(datapath_io_ex_datapathio_Forward_A),
    .io_ex_datapathio_Forward_B(datapath_io_ex_datapathio_Forward_B),
    .io_ex_datapathio_alu_b_src(datapath_io_ex_datapathio_alu_b_src),
    .io_ex_datapathio_ex_aui_pc(datapath_io_ex_datapathio_ex_aui_pc),
    .io_ex_datapathio_forward_rs2_out(datapath_io_ex_datapathio_forward_rs2_out),
    .io_ex_datapathio_alu_a_src(datapath_io_ex_datapathio_alu_a_src),
    .io_wb_datapathio_wb_alu_sum(datapath_io_wb_datapathio_wb_alu_sum),
    .io_wb_datapathio_wb_dataout(datapath_io_wb_datapathio_wb_dataout),
    .io_wb_datapathio_wb_pc_4(datapath_io_wb_datapathio_wb_pc_4),
    .io_wb_datapathio_wb_imm(datapath_io_wb_datapathio_wb_imm),
    .io_wb_datapathio_wb_aui_pc(datapath_io_wb_datapathio_wb_aui_pc),
    .io_wb_datapathio_wb_Mem_to_Reg(datapath_io_wb_datapathio_wb_Mem_to_Reg),
    .io_wb_datapathio_wb_reg_writedata(datapath_io_wb_datapathio_wb_reg_writedata)
  );
  EX_MEM_Register ex_mem_register ( // @[Tile.scala 59:31:@1080.4]
    .clock(ex_mem_register_clock),
    .reset(ex_mem_register_reset),
    .io_ex_alu_sum(ex_mem_register_io_ex_alu_sum),
    .io_ex_rs2_out(ex_mem_register_io_ex_rs2_out),
    .io_ex_rd(ex_mem_register_io_ex_rd),
    .io_ex_pc_4(ex_mem_register_io_ex_pc_4),
    .io_ex_imm(ex_mem_register_io_ex_imm),
    .io_ex_aui_pc(ex_mem_register_io_ex_aui_pc),
    .io_ex_Mem_Read(ex_mem_register_io_ex_Mem_Read),
    .io_ex_Mem_Write(ex_mem_register_io_ex_Mem_Write),
    .io_ex_Data_Size(ex_mem_register_io_ex_Data_Size),
    .io_ex_Load_Type(ex_mem_register_io_ex_Load_Type),
    .io_ex_Reg_Write(ex_mem_register_io_ex_Reg_Write),
    .io_ex_Mem_to_Reg(ex_mem_register_io_ex_Mem_to_Reg),
    .io_mem_Mem_Read(ex_mem_register_io_mem_Mem_Read),
    .io_mem_Mem_Write(ex_mem_register_io_mem_Mem_Write),
    .io_mem_Data_Size(ex_mem_register_io_mem_Data_Size),
    .io_mem_Load_Type(ex_mem_register_io_mem_Load_Type),
    .io_mem_Reg_Write(ex_mem_register_io_mem_Reg_Write),
    .io_mem_Mem_to_Reg(ex_mem_register_io_mem_Mem_to_Reg),
    .io_mem_alu_sum(ex_mem_register_io_mem_alu_sum),
    .io_mem_rs2_out(ex_mem_register_io_mem_rs2_out),
    .io_mem_rd(ex_mem_register_io_mem_rd),
    .io_mem_pc_4(ex_mem_register_io_mem_pc_4),
    .io_mem_imm(ex_mem_register_io_mem_imm),
    .io_mem_aui_pc(ex_mem_register_io_mem_aui_pc)
  );
  DataCache datacache ( // @[Tile.scala 60:31:@1083.4]
    .clock(datacache_clock),
    .io_addr(datacache_io_addr),
    .io_write_data(datacache_io_write_data),
    .io_Mem_Read(datacache_io_Mem_Read),
    .io_Mem_Write(datacache_io_Mem_Write),
    .io_Data_Size(datacache_io_Data_Size),
    .io_Load_Type(datacache_io_Load_Type),
    .io_data_out(datacache_io_data_out)
  );
  MEM_WB_Register mem_wb_register ( // @[Tile.scala 61:31:@1086.4]
    .clock(mem_wb_register_clock),
    .reset(mem_wb_register_reset),
    .io_mem_dataout(mem_wb_register_io_mem_dataout),
    .io_mem_alu_sum(mem_wb_register_io_mem_alu_sum),
    .io_mem_rd(mem_wb_register_io_mem_rd),
    .io_mem_pc_4(mem_wb_register_io_mem_pc_4),
    .io_mem_imm(mem_wb_register_io_mem_imm),
    .io_mem_aui_pc(mem_wb_register_io_mem_aui_pc),
    .io_mem_Mem_to_Reg(mem_wb_register_io_mem_Mem_to_Reg),
    .io_mem_Reg_Write(mem_wb_register_io_mem_Reg_Write),
    .io_wb_Mem_to_Reg(mem_wb_register_io_wb_Mem_to_Reg),
    .io_wb_Reg_Write(mem_wb_register_io_wb_Reg_Write),
    .io_wb_dataout(mem_wb_register_io_wb_dataout),
    .io_wb_alu_sum(mem_wb_register_io_wb_alu_sum),
    .io_wb_rd(mem_wb_register_io_wb_rd),
    .io_wb_pc_4(mem_wb_register_io_wb_pc_4),
    .io_wb_imm(mem_wb_register_io_wb_imm),
    .io_wb_aui_pc(mem_wb_register_io_wb_aui_pc)
  );
  Forward forward ( // @[Tile.scala 62:31:@1089.4]
    .io_ex_mem_Reg_Write(forward_io_ex_mem_Reg_Write),
    .io_ex_mem_rd(forward_io_ex_mem_rd),
    .io_mem_wb_Reg_Write(forward_io_mem_wb_Reg_Write),
    .io_mem_wb_rd(forward_io_mem_wb_rd),
    .io_id_ex_rs1(forward_io_id_ex_rs1),
    .io_id_ex_rs2(forward_io_id_ex_rs2),
    .io_Forward_A(forward_io_Forward_A),
    .io_Forward_B(forward_io_Forward_B)
  );
  assign io_if_pc_out = pc_io_pc_out; // @[Tile.scala 76:17:@1096.4]
  assign io_if_next_pc = datapath_io_if_datapathio_if_new_pc; // @[Tile.scala 77:17:@1097.4]
  assign io_id_rs1 = if_id_register_io_id_rs1; // @[Tile.scala 103:17:@1111.4]
  assign io_id_rs2 = if_id_register_io_id_rs2; // @[Tile.scala 104:17:@1112.4]
  assign io_id_rs1_out = regfile_io_rs1_out; // @[Tile.scala 105:17:@1113.4]
  assign io_id_rs2_out = regfile_io_rs2_out; // @[Tile.scala 106:17:@1114.4]
  assign io_ex_rs1_out = id_ex_register_io_ex_rs1_out; // @[Tile.scala 160:21:@1149.4]
  assign io_ex_rs2_out = id_ex_register_io_ex_rs2_out; // @[Tile.scala 161:21:@1150.4]
  assign io_ex_alu_sum = alu_io_Sum; // @[Tile.scala 162:21:@1151.4]
  assign io_ex_alu_conflag = alu_io_Conflag; // @[Tile.scala 163:21:@1152.4]
  assign io_ex_rd = id_ex_register_io_ex_rd; // @[Tile.scala 164:21:@1153.4]
  assign io_mem_rd = ex_mem_register_io_mem_rd; // @[Tile.scala 191:23:@1172.4]
  assign io_mem_alu_sum = ex_mem_register_io_mem_alu_sum; // @[Tile.scala 192:23:@1173.4]
  assign io_mem_writedata = ex_mem_register_io_mem_rs2_out; // @[Tile.scala 193:23:@1174.4]
  assign io_mem_dataout = datacache_io_data_out; // @[Tile.scala 194:23:@1175.4]
  assign io_wb_rd = mem_wb_register_io_wb_rd; // @[Tile.scala 216:23:@1190.4]
  assign io_wb_registerwrite = datapath_io_wb_datapathio_wb_reg_writedata; // @[Tile.scala 217:23:@1191.4]
  assign io_Forward_A = forward_io_Forward_A; // @[Tile.scala 229:16:@1198.4]
  assign io_Forward_B = forward_io_Forward_B; // @[Tile.scala 230:16:@1199.4]
  assign pc_clock = clock; // @[:@1054.4]
  assign pc_reset = reset; // @[:@1055.4]
  assign pc_io_addr_input = datapath_io_if_datapathio_if_new_pc; // @[Tile.scala 69:20:@1093.4]
  assign pc_io_pc_write = io_pc_write; // @[Tile.scala 70:20:@1094.4]
  assign instcache_clock = clock; // @[:@1057.4]
  assign instcache_io_addr = pc_io_pc_out; // @[Tile.scala 73:21:@1095.4]
  assign if_id_register_clock = clock; // @[:@1060.4]
  assign if_id_register_reset = reset; // @[:@1061.4]
  assign if_id_register_io_if_pc = pc_io_pc_out; // @[Tile.scala 84:33:@1101.4]
  assign if_id_register_io_if_inst = instcache_io_inst; // @[Tile.scala 83:33:@1100.4]
  assign if_id_register_io_if_id_write = io_if_id_write; // @[Tile.scala 81:33:@1098.4]
  assign if_id_register_io_if_flush = io_if_flush; // @[Tile.scala 82:33:@1099.4]
  assign if_id_register_io_if_pc_4 = datapath_io_if_datapathio_if_pc_4; // @[Tile.scala 85:33:@1102.4]
  assign regfile_clock = clock; // @[:@1063.4]
  assign regfile_io_rs1 = if_id_register_io_id_rs1; // @[Tile.scala 92:23:@1104.4]
  assign regfile_io_rs2 = if_id_register_io_id_rs2; // @[Tile.scala 93:23:@1105.4]
  assign regfile_io_rd = mem_wb_register_io_wb_rd; // @[Tile.scala 94:23:@1106.4]
  assign regfile_io_wdata = datapath_io_wb_datapathio_wb_reg_writedata; // @[Tile.scala 95:23:@1107.4]
  assign regfile_io_regwrite = mem_wb_register_io_wb_Reg_Write; // @[Tile.scala 96:23:@1108.4]
  assign immgen_io_inst_in = if_id_register_io_id_inst; // @[Tile.scala 99:23:@1109.4]
  assign immgen_io_imm_sel = control_io_Imm_Sel; // @[Tile.scala 100:23:@1110.4]
  assign control_io_inst = if_id_register_io_id_inst; // @[Tile.scala 89:23:@1103.4]
  assign id_ex_register_clock = clock; // @[:@1072.4]
  assign id_ex_register_reset = reset; // @[:@1073.4]
  assign id_ex_register_io_id_pc = if_id_register_io_id_pc; // @[Tile.scala 128:32:@1130.4]
  assign id_ex_register_io_id_pc_4 = if_id_register_io_id_pc_4; // @[Tile.scala 129:32:@1131.4]
  assign id_ex_register_io_id_rs1_out = regfile_io_rs1_out; // @[Tile.scala 124:32:@1126.4]
  assign id_ex_register_io_id_rs2_out = regfile_io_rs2_out; // @[Tile.scala 125:32:@1127.4]
  assign id_ex_register_io_id_imm = immgen_io_imm; // @[Tile.scala 131:32:@1133.4]
  assign id_ex_register_io_id_inst = if_id_register_io_id_inst; // @[Tile.scala 130:32:@1132.4]
  assign id_ex_register_io_id_rs1 = if_id_register_io_id_rs1; // @[Tile.scala 126:32:@1128.4]
  assign id_ex_register_io_id_rs2 = if_id_register_io_id_rs2; // @[Tile.scala 127:32:@1129.4]
  assign id_ex_register_io_ALU_Src = control_io_ALU_Src; // @[Tile.scala 111:33:@1115.4]
  assign id_ex_register_io_ALUOp = control_io_ALUOp; // @[Tile.scala 112:33:@1116.4]
  assign id_ex_register_io_Branch = control_io_Branch; // @[Tile.scala 113:33:@1117.4]
  assign id_ex_register_io_Branch_Src = control_io_Branch_Src; // @[Tile.scala 114:33:@1118.4]
  assign id_ex_register_io_Jump_Type = control_io_Jump_Type; // @[Tile.scala 115:33:@1119.4]
  assign id_ex_register_io_Mem_Read = control_io_Mem_Read; // @[Tile.scala 116:33:@1120.4]
  assign id_ex_register_io_Mem_Write = control_io_Mem_Write; // @[Tile.scala 117:33:@1121.4]
  assign id_ex_register_io_Data_Size = control_io_Data_Size; // @[Tile.scala 118:33:@1122.4]
  assign id_ex_register_io_Load_Type = control_io_Load_Type; // @[Tile.scala 119:33:@1123.4]
  assign id_ex_register_io_Reg_Write = control_io_Reg_Write; // @[Tile.scala 120:33:@1124.4]
  assign id_ex_register_io_Mem_to_Reg = control_io_Mem_to_Reg; // @[Tile.scala 121:33:@1125.4]
  assign alu_io_Src_A = datapath_io_ex_datapathio_alu_a_src; // @[Tile.scala 155:16:@1146.4]
  assign alu_io_Src_B = datapath_io_ex_datapathio_alu_b_src; // @[Tile.scala 156:16:@1147.4]
  assign alu_io_ALUOp = id_ex_register_io_ex_ALUOp; // @[Tile.scala 157:16:@1148.4]
  assign datapath_io_if_datapathio_if_pc = pc_io_pc_out; // @[Tile.scala 66:47:@1092.4]
  assign datapath_io_ex_datapathio_ex_rs1_out = id_ex_register_io_ex_rs1_out; // @[Tile.scala 137:43:@1136.4]
  assign datapath_io_ex_datapathio_ex_rs2_out = id_ex_register_io_ex_rs2_out; // @[Tile.scala 151:40:@1144.4]
  assign datapath_io_ex_datapathio_ex_imm = id_ex_register_io_ex_imm; // @[Tile.scala 136:43:@1135.4]
  assign datapath_io_ex_datapathio_ex_pc = id_ex_register_io_ex_pc; // @[Tile.scala 135:43:@1134.4]
  assign datapath_io_ex_datapathio_ex_ALU_Src = id_ex_register_io_ex_ALU_Src; // @[Tile.scala 152:40:@1145.4]
  assign datapath_io_ex_datapathio_ex_Branch = id_ex_register_io_ex_Branch; // @[Tile.scala 141:45:@1138.4]
  assign datapath_io_ex_datapathio_ex_alu_conflag = alu_io_Conflag; // @[Tile.scala 142:45:@1139.4]
  assign datapath_io_ex_datapathio_ex_Branch_Src = id_ex_register_io_ex_Branch_Src; // @[Tile.scala 138:43:@1137.4]
  assign datapath_io_ex_datapathio_ex_Jump_Type = id_ex_register_io_ex_Jump_Type; // @[Tile.scala 143:45:@1140.4]
  assign datapath_io_ex_datapathio_mem_alu_sum = ex_mem_register_io_mem_alu_sum; // @[Tile.scala 146:45:@1141.4]
  assign datapath_io_ex_datapathio_Forward_A = forward_io_Forward_A; // @[Tile.scala 147:45:@1142.4]
  assign datapath_io_ex_datapathio_Forward_B = forward_io_Forward_B; // @[Tile.scala 148:45:@1143.4]
  assign datapath_io_wb_datapathio_wb_alu_sum = mem_wb_register_io_wb_alu_sum; // @[Tile.scala 208:45:@1184.4]
  assign datapath_io_wb_datapathio_wb_dataout = mem_wb_register_io_wb_dataout; // @[Tile.scala 209:45:@1185.4]
  assign datapath_io_wb_datapathio_wb_pc_4 = mem_wb_register_io_wb_pc_4; // @[Tile.scala 210:45:@1186.4]
  assign datapath_io_wb_datapathio_wb_imm = mem_wb_register_io_wb_imm; // @[Tile.scala 211:45:@1187.4]
  assign datapath_io_wb_datapathio_wb_aui_pc = mem_wb_register_io_wb_aui_pc; // @[Tile.scala 212:45:@1188.4]
  assign datapath_io_wb_datapathio_wb_Mem_to_Reg = mem_wb_register_io_wb_Mem_to_Reg; // @[Tile.scala 213:45:@1189.4]
  assign ex_mem_register_clock = clock; // @[:@1081.4]
  assign ex_mem_register_reset = reset; // @[:@1082.4]
  assign ex_mem_register_io_ex_alu_sum = alu_io_Sum; // @[Tile.scala 168:37:@1154.4]
  assign ex_mem_register_io_ex_rs2_out = datapath_io_ex_datapathio_forward_rs2_out; // @[Tile.scala 169:37:@1155.4]
  assign ex_mem_register_io_ex_rd = id_ex_register_io_ex_rd; // @[Tile.scala 170:37:@1156.4]
  assign ex_mem_register_io_ex_pc_4 = id_ex_register_io_ex_pc_4; // @[Tile.scala 171:37:@1157.4]
  assign ex_mem_register_io_ex_imm = id_ex_register_io_ex_imm; // @[Tile.scala 172:37:@1158.4]
  assign ex_mem_register_io_ex_aui_pc = datapath_io_ex_datapathio_ex_aui_pc; // @[Tile.scala 173:37:@1159.4]
  assign ex_mem_register_io_ex_Mem_Read = id_ex_register_io_ex_Mem_Read; // @[Tile.scala 174:37:@1160.4]
  assign ex_mem_register_io_ex_Mem_Write = id_ex_register_io_ex_Mem_Write; // @[Tile.scala 175:37:@1161.4]
  assign ex_mem_register_io_ex_Data_Size = id_ex_register_io_ex_Data_Size; // @[Tile.scala 176:37:@1162.4]
  assign ex_mem_register_io_ex_Load_Type = id_ex_register_io_ex_Load_Type; // @[Tile.scala 177:37:@1163.4]
  assign ex_mem_register_io_ex_Reg_Write = id_ex_register_io_ex_Reg_Write; // @[Tile.scala 178:37:@1164.4]
  assign ex_mem_register_io_ex_Mem_to_Reg = id_ex_register_io_ex_Mem_to_Reg; // @[Tile.scala 179:37:@1165.4]
  assign datacache_clock = clock; // @[:@1084.4]
  assign datacache_io_addr = ex_mem_register_io_mem_alu_sum; // @[Tile.scala 183:27:@1166.4]
  assign datacache_io_write_data = ex_mem_register_io_mem_rs2_out; // @[Tile.scala 184:27:@1167.4]
  assign datacache_io_Mem_Read = ex_mem_register_io_mem_Mem_Read; // @[Tile.scala 185:27:@1168.4]
  assign datacache_io_Mem_Write = ex_mem_register_io_mem_Mem_Write; // @[Tile.scala 186:27:@1169.4]
  assign datacache_io_Data_Size = ex_mem_register_io_mem_Data_Size; // @[Tile.scala 187:27:@1170.4]
  assign datacache_io_Load_Type = ex_mem_register_io_mem_Load_Type; // @[Tile.scala 188:27:@1171.4]
  assign mem_wb_register_clock = clock; // @[:@1087.4]
  assign mem_wb_register_reset = reset; // @[:@1088.4]
  assign mem_wb_register_io_mem_dataout = datacache_io_data_out; // @[Tile.scala 200:39:@1178.4]
  assign mem_wb_register_io_mem_alu_sum = ex_mem_register_io_mem_alu_sum; // @[Tile.scala 201:39:@1179.4]
  assign mem_wb_register_io_mem_rd = ex_mem_register_io_mem_rd; // @[Tile.scala 202:39:@1180.4]
  assign mem_wb_register_io_mem_pc_4 = ex_mem_register_io_mem_pc_4; // @[Tile.scala 203:39:@1181.4]
  assign mem_wb_register_io_mem_imm = ex_mem_register_io_mem_imm; // @[Tile.scala 204:39:@1182.4]
  assign mem_wb_register_io_mem_aui_pc = ex_mem_register_io_mem_aui_pc; // @[Tile.scala 205:39:@1183.4]
  assign mem_wb_register_io_mem_Mem_to_Reg = ex_mem_register_io_mem_Mem_to_Reg; // @[Tile.scala 199:39:@1177.4]
  assign mem_wb_register_io_mem_Reg_Write = ex_mem_register_io_mem_Reg_Write; // @[Tile.scala 198:39:@1176.4]
  assign forward_io_ex_mem_Reg_Write = ex_mem_register_io_mem_Reg_Write; // @[Tile.scala 221:31:@1192.4]
  assign forward_io_ex_mem_rd = ex_mem_register_io_mem_rd; // @[Tile.scala 222:31:@1193.4]
  assign forward_io_mem_wb_Reg_Write = mem_wb_register_io_wb_Reg_Write; // @[Tile.scala 223:31:@1194.4]
  assign forward_io_mem_wb_rd = mem_wb_register_io_wb_rd; // @[Tile.scala 224:31:@1195.4]
  assign forward_io_id_ex_rs1 = id_ex_register_io_ex_rs1; // @[Tile.scala 225:31:@1196.4]
  assign forward_io_id_ex_rs2 = id_ex_register_io_ex_rs2; // @[Tile.scala 226:31:@1197.4]
endmodule
