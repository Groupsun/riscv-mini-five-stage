module ALU( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_Src_A, // @[:@6.4]
  input  [31:0] io_Src_B, // @[:@6.4]
  input  [3:0]  io_ALUOp, // @[:@6.4]
  output [31:0] io_Sum, // @[:@6.4]
  output        io_Zero // @[:@6.4]
);
  wire [32:0] _T_20; // @[ALU.scala 38:26:@8.4]
  wire [31:0] _T_21; // @[ALU.scala 38:26:@9.4]
  wire [32:0] _T_22; // @[ALU.scala 39:26:@10.4]
  wire [32:0] _T_23; // @[ALU.scala 39:26:@11.4]
  wire [31:0] _T_24; // @[ALU.scala 39:26:@12.4]
  wire [31:0] _T_25; // @[ALU.scala 40:26:@13.4]
  wire [31:0] _T_26; // @[ALU.scala 41:26:@14.4]
  wire  _T_27; // @[Mux.scala 46:19:@15.4]
  wire [31:0] _T_28; // @[Mux.scala 46:16:@16.4]
  wire  _T_29; // @[Mux.scala 46:19:@17.4]
  wire [31:0] _T_30; // @[Mux.scala 46:16:@18.4]
  wire  _T_31; // @[Mux.scala 46:19:@19.4]
  wire [31:0] _T_32; // @[Mux.scala 46:16:@20.4]
  wire  _T_33; // @[Mux.scala 46:19:@21.4]
  assign _T_20 = io_Src_A + io_Src_B; // @[ALU.scala 38:26:@8.4]
  assign _T_21 = io_Src_A + io_Src_B; // @[ALU.scala 38:26:@9.4]
  assign _T_22 = io_Src_A - io_Src_B; // @[ALU.scala 39:26:@10.4]
  assign _T_23 = $unsigned(_T_22); // @[ALU.scala 39:26:@11.4]
  assign _T_24 = _T_23[31:0]; // @[ALU.scala 39:26:@12.4]
  assign _T_25 = io_Src_A & io_Src_B; // @[ALU.scala 40:26:@13.4]
  assign _T_26 = io_Src_A | io_Src_B; // @[ALU.scala 41:26:@14.4]
  assign _T_27 = 4'h3 == io_ALUOp; // @[Mux.scala 46:19:@15.4]
  assign _T_28 = _T_27 ? _T_26 : io_Src_B; // @[Mux.scala 46:16:@16.4]
  assign _T_29 = 4'h2 == io_ALUOp; // @[Mux.scala 46:19:@17.4]
  assign _T_30 = _T_29 ? _T_25 : _T_28; // @[Mux.scala 46:16:@18.4]
  assign _T_31 = 4'h1 == io_ALUOp; // @[Mux.scala 46:19:@19.4]
  assign _T_32 = _T_31 ? _T_24 : _T_30; // @[Mux.scala 46:16:@20.4]
  assign _T_33 = 4'h0 == io_ALUOp; // @[Mux.scala 46:19:@21.4]
  assign io_Sum = _T_33 ? _T_21 : _T_32; // @[ALU.scala 37:10:@23.4]
  assign io_Zero = io_Src_A == io_Src_B; // @[ALU.scala 44:11:@26.4]
endmodule
